
module vgafb ( sys_clk, sys_rst, csr_a, csr_we, csr_di, csr_do, fml_adr, 
        fml_stb, fml_ack, fml_di, dcb_stb, dcb_adr, dcb_dat, dcb_hit, vga_clk, 
        vga_psave_n, vga_hsync_n, vga_vsync_n, vga_sync_n, vga_blank_n, vga_r, 
        vga_g, vga_b, vga_sda, vga_sdc );
  input [13:0] csr_a;
  input [31:0] csr_di;
  output [31:0] csr_do;
  output [25:0] fml_adr;
  input [63:0] fml_di;
  output [25:0] dcb_adr;
  input [63:0] dcb_dat;
  output [7:0] vga_r;
  output [7:0] vga_g;
  output [7:0] vga_b;
  input sys_clk, sys_rst, csr_we, fml_ack, dcb_hit, vga_clk;
  output fml_stb, dcb_stb, vga_psave_n, vga_hsync_n, vga_vsync_n, vga_sync_n,
         vga_blank_n, vga_sdc;
  inout vga_sda;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, vga_rst, baseaddress_ack, hactive,
         vactive, active, N9, generate_en, N10, N11, N12, N13, hsync_n,
         vsync_n, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25,
         N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39,
         N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53,
         N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67,
         N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81,
         N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95,
         N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107,
         N108, N109, N110, N111, N112, N113, fifo_full, pixel_valid, pixel_ack,
         N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N124,
         N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135,
         N136, N137, N138, \ctlif/N272 , \ctlif/N271 , \ctlif/N270 ,
         \ctlif/N269 , \ctlif/N268 , \ctlif/N267 , \ctlif/N266 , \ctlif/N265 ,
         \ctlif/N264 , \ctlif/N263 , \ctlif/N262 , \ctlif/N261 , \ctlif/N260 ,
         \ctlif/N259 , \ctlif/N258 , \ctlif/N257 , \ctlif/N256 , \ctlif/N255 ,
         \ctlif/N254 , \ctlif/N253 , \ctlif/N252 , \ctlif/N251 , \ctlif/N250 ,
         \ctlif/N249 , \ctlif/N248 , \ctlif/N247 , \ctlif/N246 , \ctlif/N245 ,
         \ctlif/N244 , \ctlif/N243 , \ctlif/N242 , \ctlif/N241 , \ctlif/N240 ,
         \ctlif/N239 , \ctlif/N238 , \ctlif/N237 , \ctlif/N236 , \ctlif/N235 ,
         \ctlif/N234 , \ctlif/N233 , \ctlif/N232 , \ctlif/N231 , \ctlif/N230 ,
         \ctlif/N229 , \ctlif/N228 , \ctlif/N227 , \ctlif/N226 , \ctlif/N225 ,
         \ctlif/N224 , \ctlif/N223 , \ctlif/N222 , \ctlif/N221 , \ctlif/N220 ,
         \ctlif/N219 , \ctlif/N218 , \ctlif/N217 , \ctlif/N216 , \ctlif/N215 ,
         \ctlif/N214 , \ctlif/N213 , \ctlif/N212 , \ctlif/N211 , \ctlif/N210 ,
         \ctlif/N209 , \ctlif/N208 , \ctlif/N207 , \ctlif/N206 , \ctlif/N205 ,
         \ctlif/N204 , \ctlif/N203 , \ctlif/N202 , \ctlif/N201 , \ctlif/N200 ,
         \ctlif/N199 , \ctlif/N198 , \ctlif/N197 , \ctlif/N196 , \ctlif/N195 ,
         \ctlif/N194 , \ctlif/N193 , \ctlif/N192 , \ctlif/N191 , \ctlif/N190 ,
         \ctlif/N189 , \ctlif/N188 , \ctlif/N187 , \ctlif/N186 , \ctlif/N185 ,
         \ctlif/N184 , \ctlif/N183 , \ctlif/N182 , \ctlif/N181 , \ctlif/N180 ,
         \ctlif/N179 , \ctlif/N178 , \ctlif/N177 , \ctlif/N176 , \ctlif/N175 ,
         \ctlif/N174 , \ctlif/N173 , \ctlif/N172 , \ctlif/N171 , \ctlif/N170 ,
         \ctlif/N169 , \ctlif/N168 , \ctlif/N167 , \ctlif/N166 , \ctlif/N165 ,
         \ctlif/N164 , \ctlif/N163 , \ctlif/N162 , \ctlif/N161 , \ctlif/N160 ,
         \ctlif/N159 , \ctlif/N158 , \ctlif/N157 , \ctlif/N156 , \ctlif/N155 ,
         \ctlif/N154 , \ctlif/N153 , \ctlif/N152 , \ctlif/N151 , \ctlif/N150 ,
         \ctlif/N149 , \ctlif/N148 , \ctlif/N147 , \ctlif/N146 , \ctlif/N145 ,
         \ctlif/N144 , \ctlif/N143 , \ctlif/N142 , \ctlif/N141 , \ctlif/N140 ,
         \ctlif/N139 , \ctlif/N138 , \ctlif/N137 , \ctlif/N136 , \ctlif/N135 ,
         \ctlif/N134 , \ctlif/N133 , \ctlif/N132 , \ctlif/N131 , \ctlif/N130 ,
         \ctlif/N129 , \ctlif/N128 , \ctlif/N127 , \ctlif/N126 , \ctlif/N125 ,
         \ctlif/N124 , \ctlif/N123 , \ctlif/N122 , \ctlif/N121 , \ctlif/N120 ,
         \ctlif/N119 , \ctlif/N118 , \ctlif/N117 , \ctlif/N116 , \ctlif/N115 ,
         \ctlif/N114 , \ctlif/N113 , \ctlif/N112 , \ctlif/N111 , \ctlif/N110 ,
         \ctlif/N109 , \ctlif/N108 , \ctlif/N107 , \ctlif/N106 , \ctlif/N105 ,
         \ctlif/N104 , \ctlif/N103 , \ctlif/N102 , \ctlif/N101 , \ctlif/N100 ,
         \ctlif/N99 , \ctlif/N98 , \ctlif/N97 , \ctlif/N96 , \ctlif/N95 ,
         \ctlif/N94 , \ctlif/N93 , \ctlif/N92 , \ctlif/N91 , \ctlif/N90 ,
         \ctlif/N89 , \ctlif/N88 , \ctlif/N87 , \ctlif/N86 , \ctlif/N85 ,
         \ctlif/N84 , \ctlif/N83 , \ctlif/N82 , \ctlif/N81 , \ctlif/N80 ,
         \ctlif/N79 , \ctlif/N78 , \ctlif/N77 , \ctlif/N76 , \ctlif/N75 ,
         \ctlif/N74 , \ctlif/N73 , \ctlif/N72 , \ctlif/N71 , \ctlif/N70 ,
         \ctlif/N69 , \ctlif/N68 , \ctlif/N67 , \ctlif/N66 , \ctlif/N65 ,
         \ctlif/N64 , \ctlif/N63 , \ctlif/N62 , \ctlif/N61 , \ctlif/N60 ,
         \ctlif/N59 , \ctlif/N58 , \ctlif/N57 , \ctlif/N56 , \ctlif/N55 ,
         \ctlif/N54 , \ctlif/N53 , \ctlif/N52 , \ctlif/N51 , \ctlif/N50 ,
         \ctlif/N49 , \ctlif/N48 , \ctlif/N47 , \ctlif/N46 , \ctlif/N45 ,
         \ctlif/N44 , \ctlif/N43 , \ctlif/N42 , \ctlif/N41 , \ctlif/N40 ,
         \ctlif/N39 , \ctlif/N38 , \ctlif/N37 , \ctlif/N36 , \ctlif/N35 ,
         \ctlif/N34 , \ctlif/N33 , \ctlif/N32 , \ctlif/N31 , \ctlif/N30 ,
         \ctlif/N29 , \ctlif/N28 , \ctlif/N27 , \ctlif/N26 , \ctlif/N25 ,
         \ctlif/N24 , \ctlif/sda_o , \ctlif/sda_oe , \ctlif/sda_1 ,
         \ctlif/sda_2 , \ctlif/N23 , \ctlif/N22 , \ctlif/N21 , \ctlif/N20 ,
         \ctlif/N19 , \ctlif/N18 , \ctlif/N17 , \ctlif/N16 , \ctlif/N15 ,
         \ctlif/N14 , \ctlif/N13 , \ctlif/N12 , \ctlif/N11 , \ctlif/N10 ,
         \ctlif/N9 , \ctlif/N8 , \ctlif/N7 , \ctlif/N6 , \ctlif/N5 ,
         \ctlif/N4 , \ctlif/N3 , \ctlif/N2 , \ctlif/N1 , \ctlif/N0 ,
         \pixelfeed/N266 , \pixelfeed/N265 , \pixelfeed/N264 ,
         \pixelfeed/N263 , \pixelfeed/N262 , \pixelfeed/N261 ,
         \pixelfeed/N260 , \pixelfeed/N259 , \pixelfeed/N258 ,
         \pixelfeed/N257 , \pixelfeed/N256 , \pixelfeed/N255 ,
         \pixelfeed/N254 , \pixelfeed/N253 , \pixelfeed/N252 ,
         \pixelfeed/N251 , \pixelfeed/N250 , \pixelfeed/N249 ,
         \pixelfeed/N248 , \pixelfeed/N247 , \pixelfeed/N246 ,
         \pixelfeed/N245 , \pixelfeed/N244 , \pixelfeed/N243 ,
         \pixelfeed/N242 , \pixelfeed/N241 , \pixelfeed/N240 ,
         \pixelfeed/N239 , \pixelfeed/N238 , \pixelfeed/N237 ,
         \pixelfeed/N236 , \pixelfeed/N235 , \pixelfeed/N234 ,
         \pixelfeed/N233 , \pixelfeed/N232 , \pixelfeed/N231 ,
         \pixelfeed/N230 , \pixelfeed/N229 , \pixelfeed/N228 ,
         \pixelfeed/N227 , \pixelfeed/N226 , \pixelfeed/N225 ,
         \pixelfeed/N224 , \pixelfeed/N223 , \pixelfeed/N222 ,
         \pixelfeed/N221 , \pixelfeed/N220 , \pixelfeed/N219 ,
         \pixelfeed/N218 , \pixelfeed/N217 , \pixelfeed/N216 ,
         \pixelfeed/N215 , \pixelfeed/N214 , \pixelfeed/N213 ,
         \pixelfeed/N212 , \pixelfeed/N211 , \pixelfeed/N210 ,
         \pixelfeed/N209 , \pixelfeed/N208 , \pixelfeed/N207 ,
         \pixelfeed/N206 , \pixelfeed/N205 , \pixelfeed/N204 ,
         \pixelfeed/N203 , \pixelfeed/N202 , \pixelfeed/N201 ,
         \pixelfeed/N200 , \pixelfeed/N199 , \pixelfeed/N198 ,
         \pixelfeed/N197 , \pixelfeed/N196 , \pixelfeed/N195 ,
         \pixelfeed/N194 , \pixelfeed/N193 , \pixelfeed/N192 ,
         \pixelfeed/N191 , \pixelfeed/N190 , \pixelfeed/N189 ,
         \pixelfeed/N188 , \pixelfeed/N187 , \pixelfeed/N186 ,
         \pixelfeed/N185 , \pixelfeed/N184 , \pixelfeed/N183 ,
         \pixelfeed/N182 , \pixelfeed/N181 , \pixelfeed/N180 ,
         \pixelfeed/N179 , \pixelfeed/N178 , \pixelfeed/N177 ,
         \pixelfeed/N176 , \pixelfeed/N175 , \pixelfeed/N174 ,
         \pixelfeed/N173 , \pixelfeed/N172 , \pixelfeed/N171 ,
         \pixelfeed/N170 , \pixelfeed/N169 , \pixelfeed/N168 ,
         \pixelfeed/N167 , \pixelfeed/N166 , \pixelfeed/N165 ,
         \pixelfeed/N164 , \pixelfeed/N163 , \pixelfeed/N162 ,
         \pixelfeed/N161 , \pixelfeed/N160 , \pixelfeed/N159 ,
         \pixelfeed/N158 , \pixelfeed/N157 , \pixelfeed/N156 ,
         \pixelfeed/ignore , \pixelfeed/ignore_clear , \pixelfeed/N155 ,
         \pixelfeed/N154 , \pixelfeed/N153 , \pixelfeed/N152 ,
         \pixelfeed/state[0] , \pixelfeed/state[1] , \pixelfeed/state[2] ,
         \pixelfeed/state[3] , \pixelfeed/N151 , \pixelfeed/N150 ,
         \pixelfeed/N149 , \pixelfeed/N148 , \pixelfeed/N147 ,
         \pixelfeed/N146 , \pixelfeed/N145 , \pixelfeed/N144 ,
         \pixelfeed/N143 , \pixelfeed/N142 , \pixelfeed/N141 ,
         \pixelfeed/N140 , \pixelfeed/N139 , \pixelfeed/N138 ,
         \pixelfeed/N137 , \pixelfeed/N136 , \pixelfeed/N135 ,
         \pixelfeed/N134 , \pixelfeed/N133 , \pixelfeed/N132 ,
         \pixelfeed/N131 , \pixelfeed/N130 , \pixelfeed/N129 ,
         \pixelfeed/N128 , \pixelfeed/N127 , \pixelfeed/N126 ,
         \pixelfeed/N125 , \pixelfeed/N124 , \pixelfeed/N123 ,
         \pixelfeed/N122 , \pixelfeed/N121 , \pixelfeed/N120 ,
         \pixelfeed/N119 , \pixelfeed/N118 , \pixelfeed/N117 ,
         \pixelfeed/N116 , \pixelfeed/N115 , \pixelfeed/N114 ,
         \pixelfeed/N113 , \pixelfeed/N112 , \pixelfeed/N111 ,
         \pixelfeed/N110 , \pixelfeed/N109 , \pixelfeed/N108 ,
         \pixelfeed/N107 , \pixelfeed/N106 , \pixelfeed/N105 ,
         \pixelfeed/N104 , \pixelfeed/N103 , \pixelfeed/N102 ,
         \pixelfeed/N101 , \pixelfeed/N100 , \pixelfeed/N99 , \pixelfeed/N98 ,
         \pixelfeed/N97 , \pixelfeed/N96 , \pixelfeed/N95 , \pixelfeed/N94 ,
         \pixelfeed/N93 , \pixelfeed/N92 , \pixelfeed/N91 , \pixelfeed/N90 ,
         \pixelfeed/N89 , \pixelfeed/N88 , \pixelfeed/N87 , \pixelfeed/N86 ,
         \pixelfeed/N85 , \pixelfeed/N84 , \pixelfeed/N83 , \pixelfeed/N82 ,
         \pixelfeed/N81 , \pixelfeed/N80 , \pixelfeed/N79 , \pixelfeed/N78 ,
         \pixelfeed/N77 , \pixelfeed/N76 , \pixelfeed/N75 , \pixelfeed/N74 ,
         \pixelfeed/N73 , \pixelfeed/N72 , \pixelfeed/N71 , \pixelfeed/N70 ,
         \pixelfeed/N69 , \pixelfeed/N68 , \pixelfeed/N67 , \pixelfeed/N66 ,
         \pixelfeed/N65 , \pixelfeed/N64 , \pixelfeed/N63 , \pixelfeed/N62 ,
         \pixelfeed/N61 , \pixelfeed/N60 , \pixelfeed/N59 , \pixelfeed/N58 ,
         \pixelfeed/N57 , \pixelfeed/N56 , \pixelfeed/N55 , \pixelfeed/N54 ,
         \pixelfeed/N53 , \pixelfeed/N52 , \pixelfeed/N51 , \pixelfeed/N50 ,
         \pixelfeed/N49 , \pixelfeed/N48 , \pixelfeed/N47 , \pixelfeed/N46 ,
         \pixelfeed/N45 , \pixelfeed/N44 , \pixelfeed/N43 , \pixelfeed/N42 ,
         \pixelfeed/N41 , \pixelfeed/N40 , \pixelfeed/N39 , \pixelfeed/N38 ,
         \pixelfeed/N37 , \pixelfeed/sof , \pixelfeed/N36 ,
         \pixelfeed/bcounter[0] , \pixelfeed/bcounter[1] ,
         \pixelfeed/bcounter[2] , \pixelfeed/bcounter[3] ,
         \pixelfeed/bcounter[4] , \pixelfeed/bcounter[5] ,
         \pixelfeed/bcounter[6] , \pixelfeed/bcounter[7] ,
         \pixelfeed/bcounter[8] , \pixelfeed/bcounter[9] ,
         \pixelfeed/bcounter[10] , \pixelfeed/bcounter[11] ,
         \pixelfeed/bcounter[12] , \pixelfeed/bcounter[13] ,
         \pixelfeed/bcounter[14] , \pixelfeed/bcounter[15] ,
         \pixelfeed/bcounter[16] , \pixelfeed/bcounter[17] , \pixelfeed/N35 ,
         \pixelfeed/fifo_source_cache , \pixelfeed/n_0_net__0_ ,
         \pixelfeed/n_0_net__1_ , \pixelfeed/n_0_net__2_ ,
         \pixelfeed/n_0_net__3_ , \pixelfeed/n_0_net__4_ ,
         \pixelfeed/n_0_net__5_ , \pixelfeed/n_0_net__6_ ,
         \pixelfeed/n_0_net__7_ , \pixelfeed/n_0_net__8_ ,
         \pixelfeed/n_0_net__9_ , \pixelfeed/n_0_net__10_ ,
         \pixelfeed/n_0_net__11_ , \pixelfeed/n_0_net__12_ ,
         \pixelfeed/n_0_net__13_ , \pixelfeed/n_0_net__14_ ,
         \pixelfeed/n_0_net__15_ , \pixelfeed/n_0_net__16_ ,
         \pixelfeed/n_0_net__17_ , \pixelfeed/n_0_net__18_ ,
         \pixelfeed/n_0_net__19_ , \pixelfeed/n_0_net__20_ ,
         \pixelfeed/n_0_net__21_ , \pixelfeed/n_0_net__22_ ,
         \pixelfeed/n_0_net__23_ , \pixelfeed/n_0_net__24_ ,
         \pixelfeed/n_0_net__25_ , \pixelfeed/n_0_net__26_ ,
         \pixelfeed/n_0_net__27_ , \pixelfeed/n_0_net__28_ ,
         \pixelfeed/n_0_net__29_ , \pixelfeed/n_0_net__30_ ,
         \pixelfeed/n_0_net__31_ , \pixelfeed/n_0_net__32_ ,
         \pixelfeed/n_0_net__33_ , \pixelfeed/n_0_net__34_ ,
         \pixelfeed/n_0_net__35_ , \pixelfeed/n_0_net__36_ ,
         \pixelfeed/n_0_net__37_ , \pixelfeed/n_0_net__38_ ,
         \pixelfeed/n_0_net__39_ , \pixelfeed/n_0_net__40_ ,
         \pixelfeed/n_0_net__41_ , \pixelfeed/n_0_net__42_ ,
         \pixelfeed/n_0_net__43_ , \pixelfeed/n_0_net__44_ ,
         \pixelfeed/n_0_net__45_ , \pixelfeed/n_0_net__46_ ,
         \pixelfeed/n_0_net__47_ , \pixelfeed/n_0_net__48_ ,
         \pixelfeed/n_0_net__49_ , \pixelfeed/n_0_net__50_ ,
         \pixelfeed/n_0_net__51_ , \pixelfeed/n_0_net__52_ ,
         \pixelfeed/n_0_net__53_ , \pixelfeed/n_0_net__54_ ,
         \pixelfeed/n_0_net__55_ , \pixelfeed/n_0_net__56_ ,
         \pixelfeed/n_0_net__57_ , \pixelfeed/n_0_net__58_ ,
         \pixelfeed/n_0_net__59_ , \pixelfeed/n_0_net__60_ ,
         \pixelfeed/n_0_net__61_ , \pixelfeed/n_0_net__62_ ,
         \pixelfeed/n_0_net__63_ , \pixelfeed/fifo_stb , \pixelfeed/N34 ,
         \pixelfeed/N33 , \pixelfeed/N32 , \pixelfeed/N31 , \pixelfeed/N30 ,
         \pixelfeed/N29 , \pixelfeed/N28 , \pixelfeed/N27 , \pixelfeed/N26 ,
         \pixelfeed/N25 , \pixelfeed/N24 , \pixelfeed/N23 , \pixelfeed/N22 ,
         \pixelfeed/N21 , \pixelfeed/N20 , \pixelfeed/N19 , \pixelfeed/N18 ,
         \pixelfeed/N17 , \pixelfeed/N16 , \pixelfeed/N15 , \pixelfeed/N14 ,
         \pixelfeed/N13 , \pixelfeed/N12 , \pixelfeed/N11 , \pixelfeed/N10 ,
         \pixelfeed/N9 , \pixelfeed/N8 , \pixelfeed/N7 , \pixelfeed/N6 ,
         \pixelfeed/N5 , \pixelfeed/N4 , \pixelfeed/N3 , \pixelfeed/N2 ,
         \pixelfeed/N1 , \pixelfeed/N0 , \pixelfeed/fifo64to16/N95 ,
         \pixelfeed/fifo64to16/N94 , \pixelfeed/fifo64to16/N93 ,
         \pixelfeed/fifo64to16/N92 , \pixelfeed/fifo64to16/N91 ,
         \pixelfeed/fifo64to16/N90 , \pixelfeed/fifo64to16/N89 ,
         \pixelfeed/fifo64to16/N88 , \pixelfeed/fifo64to16/N87 ,
         \pixelfeed/fifo64to16/N86 , \pixelfeed/fifo64to16/N85 ,
         \pixelfeed/fifo64to16/N84 , \pixelfeed/fifo64to16/N83 ,
         \pixelfeed/fifo64to16/N82 , \pixelfeed/fifo64to16/N81 ,
         \pixelfeed/fifo64to16/N80 , \pixelfeed/fifo64to16/N79 ,
         \pixelfeed/fifo64to16/N78 , \pixelfeed/fifo64to16/N77 ,
         \pixelfeed/fifo64to16/N76 , \pixelfeed/fifo64to16/N75 ,
         \pixelfeed/fifo64to16/N74 , \pixelfeed/fifo64to16/N73 ,
         \pixelfeed/fifo64to16/N72 , \pixelfeed/fifo64to16/N71 ,
         \pixelfeed/fifo64to16/N70 , \pixelfeed/fifo64to16/N69 ,
         \pixelfeed/fifo64to16/N68 , \pixelfeed/fifo64to16/N67 ,
         \pixelfeed/fifo64to16/N66 , \pixelfeed/fifo64to16/N65 ,
         \pixelfeed/fifo64to16/N64 , \pixelfeed/fifo64to16/N63 ,
         \pixelfeed/fifo64to16/N62 , \pixelfeed/fifo64to16/N61 ,
         \pixelfeed/fifo64to16/N60 , \pixelfeed/fifo64to16/N59 ,
         \pixelfeed/fifo64to16/N58 , \pixelfeed/fifo64to16/N57 ,
         \pixelfeed/fifo64to16/N56 , \pixelfeed/fifo64to16/N55 ,
         \pixelfeed/fifo64to16/N54 , \pixelfeed/fifo64to16/N53 ,
         \pixelfeed/fifo64to16/N52 , \pixelfeed/fifo64to16/N51 ,
         \pixelfeed/fifo64to16/N50 , \pixelfeed/fifo64to16/N49 ,
         \pixelfeed/fifo64to16/N48 , \pixelfeed/fifo64to16/N47 ,
         \pixelfeed/fifo64to16/N46 , \pixelfeed/fifo64to16/N45 ,
         \pixelfeed/fifo64to16/N44 , \pixelfeed/fifo64to16/N43 ,
         \pixelfeed/fifo64to16/N42 , \pixelfeed/fifo64to16/N41 ,
         \pixelfeed/fifo64to16/N40 , \pixelfeed/fifo64to16/N39 ,
         \pixelfeed/fifo64to16/N38 , \pixelfeed/fifo64to16/N37 ,
         \pixelfeed/fifo64to16/N36 , \pixelfeed/fifo64to16/N35 ,
         \pixelfeed/fifo64to16/N34 , \pixelfeed/fifo64to16/N33 ,
         \pixelfeed/fifo64to16/N32 , \pixelfeed/fifo64to16/N31 ,
         \pixelfeed/fifo64to16/N30 , \pixelfeed/fifo64to16/N29 ,
         \pixelfeed/fifo64to16/N28 , \pixelfeed/fifo64to16/N27 ,
         \pixelfeed/fifo64to16/N26 , \pixelfeed/fifo64to16/N25 ,
         \pixelfeed/fifo64to16/level[0] , \pixelfeed/fifo64to16/level[1] ,
         \pixelfeed/fifo64to16/level[2] , \pixelfeed/fifo64to16/level[3] ,
         \pixelfeed/fifo64to16/level[4] , \pixelfeed/fifo64to16/N24 ,
         \pixelfeed/fifo64to16/produce[0] , \pixelfeed/fifo64to16/produce[1] ,
         \pixelfeed/fifo64to16/N23 , \pixelfeed/fifo64to16/N22 ,
         \pixelfeed/fifo64to16/N21 , \pixelfeed/fifo64to16/N20 ,
         \pixelfeed/fifo64to16/N19 , \pixelfeed/fifo64to16/N18 ,
         \pixelfeed/fifo64to16/N17 , \pixelfeed/fifo64to16/N16 ,
         \pixelfeed/fifo64to16/consume[0] , \pixelfeed/fifo64to16/consume[1] ,
         \pixelfeed/fifo64to16/consume[2] , \pixelfeed/fifo64to16/consume[3] ,
         \pixelfeed/fifo64to16/N15 , \pixelfeed/fifo64to16/N14 ,
         \pixelfeed/fifo64to16/N13 , \pixelfeed/fifo64to16/N12 ,
         \pixelfeed/fifo64to16/N11 , \pixelfeed/fifo64to16/N10 ,
         \pixelfeed/fifo64to16/N9 , \pixelfeed/fifo64to16/N8 ,
         \pixelfeed/fifo64to16/N7 , \pixelfeed/fifo64to16/N6 ,
         \pixelfeed/fifo64to16/N5 , \pixelfeed/fifo64to16/N4 ,
         \pixelfeed/fifo64to16/N3 , \pixelfeed/fifo64to16/N2 ,
         \pixelfeed/fifo64to16/N1 , \pixelfeed/fifo64to16/N0 ;
  wire   [10:0] hres;
  wire   [10:0] hsync_start;
  wire   [10:0] hsync_end;
  wire   [10:0] hscan;
  wire   [10:0] vres;
  wire   [10:0] vsync_start;
  wire   [10:0] vsync_end;
  wire   [10:0] vscan;
  wire   [25:0] baseaddress;
  wire   [17:0] nbursts;
  wire   [15:0] pixel;
  wire   [15:0] pixel_fb;
  wire   [10:0] hcounter;
  wire   [10:0] vcounter;
  wire   [17:0] fifo_do;
  wire   [25:0] \ctlif/baseaddress_act ;
  wire   [3:0] \pixelfeed/next_state ;
  wire   [63:0] \pixelfeed/fifo64to16/do64 ;
  wire   [255:0] \pixelfeed/fifo64to16/storage ;
  assign vga_blank_n = 1'b1;
  assign vga_psave_n = 1'b1;
  assign vga_sync_n = 1'b0;
  assign dcb_adr[25] = fml_adr[25];
  assign dcb_adr[24] = fml_adr[24];
  assign dcb_adr[23] = fml_adr[23];
  assign dcb_adr[22] = fml_adr[22];
  assign dcb_adr[21] = fml_adr[21];
  assign dcb_adr[20] = fml_adr[20];
  assign dcb_adr[19] = fml_adr[19];
  assign dcb_adr[18] = fml_adr[18];
  assign dcb_adr[17] = fml_adr[17];
  assign dcb_adr[16] = fml_adr[16];
  assign dcb_adr[15] = fml_adr[15];
  assign dcb_adr[14] = fml_adr[14];
  assign dcb_adr[13] = fml_adr[13];
  assign dcb_adr[12] = fml_adr[12];
  assign dcb_adr[11] = fml_adr[11];
  assign dcb_adr[10] = fml_adr[10];
  assign dcb_adr[9] = fml_adr[9];
  assign dcb_adr[8] = fml_adr[8];
  assign dcb_adr[7] = fml_adr[7];
  assign dcb_adr[6] = fml_adr[6];
  assign dcb_adr[5] = fml_adr[5];
  assign dcb_adr[2] = 1'b0;
  assign dcb_adr[1] = 1'b0;
  assign dcb_adr[0] = 1'b0;

  EQ_UNS_OP eq_148 ( .A(hcounter), .B(hres), .Z(N26) );
  EQ_UNS_OP eq_149 ( .A(hcounter), .B(hsync_start), .Z(N30) );
  EQ_UNS_OP eq_150 ( .A(hcounter), .B(hsync_end), .Z(N31) );
  EQ_UNS_OP eq_151 ( .A(hcounter), .B(hscan), .Z(N34) );
  EQ_UNS_OP eq_153 ( .A(vcounter), .B(vscan), .Z(N37) );
  EQ_UNS_OP eq_160 ( .A(vcounter), .B(vres), .Z(N72) );
  EQ_UNS_OP eq_161 ( .A(vcounter), .B(vsync_start), .Z(N76) );
  EQ_UNS_OP eq_162 ( .A(vcounter), .B(vsync_end), .Z(N77) );
  \**SEQGEN**  hactive_reg ( .clear(1'b0), .preset(1'b0), .next_state(N105), 
        .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(hactive), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N104) );
  \**SEQGEN**  vsync_n_reg ( .clear(1'b0), .preset(1'b0), .next_state(N111), 
        .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(vsync_n), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N110) );
  \**SEQGEN**  vactive_reg ( .clear(1'b0), .preset(1'b0), .next_state(N109), 
        .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(vactive), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N108) );
  \**SEQGEN**  vcounter_reg_10_ ( .clear(1'b0), .preset(1'b0), .next_state(
        N102), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vcounter[10]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N103) );
  \**SEQGEN**  vcounter_reg_9_ ( .clear(1'b0), .preset(1'b0), .next_state(N101), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(vcounter[9]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N103) );
  \**SEQGEN**  vcounter_reg_8_ ( .clear(1'b0), .preset(1'b0), .next_state(N100), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(vcounter[8]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N103) );
  \**SEQGEN**  vcounter_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(N99), 
        .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(vcounter[7]), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N103) );
  \**SEQGEN**  vcounter_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(N98), 
        .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(vcounter[6]), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N103) );
  \**SEQGEN**  vcounter_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(N97), 
        .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(vcounter[5]), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N103) );
  \**SEQGEN**  vcounter_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(N96), 
        .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(vcounter[4]), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N103) );
  \**SEQGEN**  vcounter_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(N95), 
        .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(vcounter[3]), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N103) );
  \**SEQGEN**  vcounter_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(N94), 
        .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(vcounter[2]), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N103) );
  \**SEQGEN**  vcounter_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(N93), 
        .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(vcounter[1]), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N103) );
  \**SEQGEN**  vcounter_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(N92), 
        .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(vcounter[0]), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N103) );
  \**SEQGEN**  hsync_n_reg ( .clear(1'b0), .preset(1'b0), .next_state(N107), 
        .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(hsync_n), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N106) );
  \**SEQGEN**  hcounter_reg_10_ ( .clear(1'b0), .preset(1'b0), .next_state(N90), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(hcounter[10]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N91) );
  \**SEQGEN**  hcounter_reg_9_ ( .clear(1'b0), .preset(1'b0), .next_state(N89), 
        .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(hcounter[9]), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N91) );
  \**SEQGEN**  hcounter_reg_8_ ( .clear(1'b0), .preset(1'b0), .next_state(N88), 
        .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(hcounter[8]), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N91) );
  \**SEQGEN**  hcounter_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(N87), 
        .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(hcounter[7]), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N91) );
  \**SEQGEN**  hcounter_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(N86), 
        .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(hcounter[6]), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N91) );
  \**SEQGEN**  hcounter_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(N85), 
        .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(hcounter[5]), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N91) );
  \**SEQGEN**  hcounter_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(N84), 
        .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(hcounter[4]), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N91) );
  \**SEQGEN**  hcounter_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(N83), 
        .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(hcounter[3]), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N91) );
  \**SEQGEN**  hcounter_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(N82), 
        .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(hcounter[2]), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N91) );
  \**SEQGEN**  hcounter_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(N81), 
        .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(hcounter[1]), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N91) );
  \**SEQGEN**  hcounter_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(N80), 
        .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(hcounter[0]), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N91) );
  asfifo fifo ( .data_out(fifo_do), .read_en(1'b1), .clk_read(vga_clk), 
        .data_in({vsync_n, hsync_n, pixel}), .full(fifo_full), .write_en(
        generate_en), .clk_write(sys_clk), .rst(vga_rst) );
  \**SEQGEN**  vga_b_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[4]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_b[7]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_b_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[3]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_b[6]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_b_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[2]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_b[5]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_b_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[1]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_b[4]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_b_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[0]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_b[3]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_b_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[4]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_b[2]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_b_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[3]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_b[1]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_b_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[2]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_b[0]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_vsync_n_reg ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[17]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_vsync_n), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_hsync_n_reg ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[16]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_hsync_n), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_r_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[15]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_r[7]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_r_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[14]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_r[6]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_r_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[13]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_r[5]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_r_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[12]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_r[4]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_r_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[11]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_r[3]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_r_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[15]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_r[2]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_r_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[14]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_r[1]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_r_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[13]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_r[0]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_g_reg_7_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[10]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_g[7]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_g_reg_6_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[9]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_g[6]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_g_reg_5_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[8]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_g[5]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_g_reg_4_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[7]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_g[4]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_g_reg_3_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[6]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_g[3]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_g_reg_2_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[5]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_g[2]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_g_reg_1_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[10]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_g[1]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  vga_g_reg_0_ ( .clear(1'b0), .preset(1'b0), .next_state(
        fifo_do[9]), .clocked_on(vga_clk), .data_in(1'b0), .enable(1'b0), .Q(
        vga_g[0]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  GTECH_OR2 C226 ( .A(hcounter[9]), .B(hcounter[10]), .Z(N114) );
  GTECH_OR2 C227 ( .A(hcounter[8]), .B(N114), .Z(N115) );
  GTECH_OR2 C228 ( .A(hcounter[7]), .B(N115), .Z(N116) );
  GTECH_OR2 C229 ( .A(hcounter[6]), .B(N116), .Z(N117) );
  GTECH_OR2 C230 ( .A(hcounter[5]), .B(N117), .Z(N118) );
  GTECH_OR2 C231 ( .A(hcounter[4]), .B(N118), .Z(N119) );
  GTECH_OR2 C232 ( .A(hcounter[3]), .B(N119), .Z(N120) );
  GTECH_OR2 C233 ( .A(hcounter[2]), .B(N120), .Z(N121) );
  GTECH_OR2 C234 ( .A(hcounter[1]), .B(N121), .Z(N122) );
  GTECH_OR2 C235 ( .A(hcounter[0]), .B(N122), .Z(N123) );
  GTECH_NOT I_0 ( .A(N123), .Z(N124) );
  GTECH_OR2 C237 ( .A(vcounter[9]), .B(vcounter[10]), .Z(N125) );
  GTECH_OR2 C238 ( .A(vcounter[8]), .B(N125), .Z(N126) );
  GTECH_OR2 C239 ( .A(vcounter[7]), .B(N126), .Z(N127) );
  GTECH_OR2 C240 ( .A(vcounter[6]), .B(N127), .Z(N128) );
  GTECH_OR2 C241 ( .A(vcounter[5]), .B(N128), .Z(N129) );
  GTECH_OR2 C242 ( .A(vcounter[4]), .B(N129), .Z(N130) );
  GTECH_OR2 C243 ( .A(vcounter[3]), .B(N130), .Z(N131) );
  GTECH_OR2 C244 ( .A(vcounter[2]), .B(N131), .Z(N132) );
  GTECH_OR2 C245 ( .A(vcounter[1]), .B(N132), .Z(N133) );
  GTECH_OR2 C246 ( .A(vcounter[0]), .B(N133), .Z(N134) );
  GTECH_NOT I_1 ( .A(N134), .Z(N135) );
  GTECH_OR2 C248 ( .A(N10), .B(N113), .Z(N91) );
  ADD_UNS_OP add_145 ( .A(hcounter), .B(1'b1), .Z({N25, N24, N23, N22, N21, 
        N20, N19, N18, N17, N16, N15}) );
  ADD_UNS_OP add_156 ( .A(vcounter), .B(1'b1), .Z({N49, N48, N47, N46, N45, 
        N44, N43, N42, N41, N40, N39}) );
  SELECT_OP C272 ( .DATA1(pixel_fb), .DATA2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CONTROL1(N0), .CONTROL2(N1), .Z(pixel) );
  GTECH_BUF B_0 ( .A(active), .Z(N0) );
  GTECH_BUF B_1 ( .A(N9), .Z(N1) );
  SELECT_OP C273 ( .DATA1(1'b1), .DATA2(N124), .CONTROL1(N2), .CONTROL2(N27), 
        .Z(N28) );
  GTECH_BUF B_2 ( .A(N26), .Z(N2) );
  GTECH_NOT I_2 ( .A(N26), .Z(N29) );
  SELECT_OP C275 ( .DATA1(1'b1), .DATA2(N30), .CONTROL1(N3), .CONTROL2(N32), 
        .Z(N33) );
  GTECH_BUF B_3 ( .A(N31), .Z(N3) );
  SELECT_OP C276 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .DATA2({N49, N48, N47, N46, N45, N44, N43, N42, 
        N41, N40, N39}), .CONTROL1(N4), .CONTROL2(N38), .Z({N60, N59, N58, N57, 
        N56, N55, N54, N53, N52, N51, N50}) );
  GTECH_BUF B_4 ( .A(N37), .Z(N4) );
  SELECT_OP C277 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .DATA2({N25, N24, N23, N22, N21, N20, N19, N18, 
        N17, N16, N15}), .CONTROL1(N5), .CONTROL2(N35), .Z({N71, N70, N69, N68, 
        N67, N66, N65, N64, N63, N62, N61}) );
  GTECH_BUF B_5 ( .A(N34), .Z(N5) );
  SELECT_OP C278 ( .DATA1(1'b1), .DATA2(N135), .CONTROL1(N6), .CONTROL2(N73), 
        .Z(N74) );
  GTECH_BUF B_6 ( .A(N72), .Z(N6) );
  GTECH_NOT I_3 ( .A(N72), .Z(N75) );
  SELECT_OP C280 ( .DATA1(1'b1), .DATA2(N76), .CONTROL1(N7), .CONTROL2(N78), 
        .Z(N79) );
  GTECH_BUF B_7 ( .A(N77), .Z(N7) );
  SELECT_OP C281 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .DATA2({N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61}), .CONTROL1(N8), .CONTROL2(N113), .Z({N90, N89, N88, 
        N87, N86, N85, N84, N83, N82, N81, N80}) );
  GTECH_BUF B_8 ( .A(N10), .Z(N8) );
  SELECT_OP C282 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .DATA2({N60, N59, N58, N57, N56, N55, N54, N53, 
        N52, N51, N50}), .CONTROL1(N8), .CONTROL2(N113), .Z({N102, N101, N100, 
        N99, N98, N97, N96, N95, N94, N93, N92}) );
  SELECT_OP C283 ( .DATA1(1'b1), .DATA2(N34), .DATA3(1'b0), .CONTROL1(N8), 
        .CONTROL2(N113), .CONTROL3(N13), .Z(N103) );
  SELECT_OP C284 ( .DATA1(1'b1), .DATA2(N28), .DATA3(1'b0), .CONTROL1(N8), 
        .CONTROL2(N113), .CONTROL3(N13), .Z(N104) );
  SELECT_OP C285 ( .DATA1(1'b0), .DATA2(N29), .CONTROL1(N8), .CONTROL2(N113), 
        .Z(N105) );
  SELECT_OP C286 ( .DATA1(1'b1), .DATA2(N33), .DATA3(1'b0), .CONTROL1(N8), 
        .CONTROL2(N113), .CONTROL3(N13), .Z(N106) );
  SELECT_OP C287 ( .DATA1(1'b1), .DATA2(N31), .CONTROL1(N8), .CONTROL2(N113), 
        .Z(N107) );
  SELECT_OP C288 ( .DATA1(1'b1), .DATA2(N74), .DATA3(1'b0), .CONTROL1(N8), 
        .CONTROL2(N113), .CONTROL3(N13), .Z(N108) );
  SELECT_OP C289 ( .DATA1(1'b0), .DATA2(N75), .CONTROL1(N8), .CONTROL2(N113), 
        .Z(N109) );
  SELECT_OP C290 ( .DATA1(1'b1), .DATA2(N79), .DATA3(1'b0), .CONTROL1(N8), 
        .CONTROL2(N113), .CONTROL3(N13), .Z(N110) );
  SELECT_OP C291 ( .DATA1(1'b1), .DATA2(N77), .CONTROL1(N8), .CONTROL2(N113), 
        .Z(N111) );
  GTECH_AND2 C294 ( .A(hactive), .B(vactive), .Z(active) );
  GTECH_NOT I_4 ( .A(active), .Z(N9) );
  GTECH_BUF B_9 ( .A(vga_rst), .Z(N10) );
  GTECH_BUF B_10 ( .A(generate_en), .Z(N11) );
  GTECH_OR2 C300 ( .A(N11), .B(N10), .Z(N12) );
  GTECH_NOT I_5 ( .A(N12), .Z(N13) );
  GTECH_BUF B_11 ( .A(N113), .Z(N14) );
  GTECH_NOT I_6 ( .A(N26), .Z(N27) );
  GTECH_NOT I_7 ( .A(N31), .Z(N32) );
  GTECH_NOT I_8 ( .A(N34), .Z(N35) );
  GTECH_AND2 C311 ( .A(N14), .B(N34), .Z(N36) );
  GTECH_NOT I_9 ( .A(N37), .Z(N38) );
  GTECH_AND2 C314 ( .A(N36), .B(N38), .Z() );
  GTECH_NOT I_10 ( .A(N72), .Z(N73) );
  GTECH_NOT I_11 ( .A(N77), .Z(N78) );
  GTECH_NOT I_12 ( .A(N10), .Z(N112) );
  GTECH_AND2 C324 ( .A(N11), .B(N112), .Z(N113) );
  GTECH_AND2 C325 ( .A(N14), .B(N112), .Z() );
  GTECH_AND2 C326 ( .A(N136), .B(N137), .Z(generate_en) );
  GTECH_NOT I_13 ( .A(fifo_full), .Z(N136) );
  GTECH_OR2 C328 ( .A(N9), .B(pixel_valid), .Z(N137) );
  GTECH_AND2 C330 ( .A(N138), .B(pixel_valid), .Z(pixel_ack) );
  GTECH_AND2 C331 ( .A(N136), .B(active), .Z(N138) );
  GTECH_NOT \ctlif/I_22  ( .A(\ctlif/N118 ), .Z(\ctlif/N119 ) );
  GTECH_OR2 \ctlif/C1644  ( .A(\ctlif/N106 ), .B(\ctlif/N117 ), .Z(
        \ctlif/N118 ) );
  GTECH_OR2 \ctlif/C1643  ( .A(\ctlif/N100 ), .B(\ctlif/N116 ), .Z(
        \ctlif/N117 ) );
  GTECH_OR2 \ctlif/C1642  ( .A(\ctlif/N94 ), .B(\ctlif/N115 ), .Z(\ctlif/N116 ) );
  GTECH_OR2 \ctlif/C1641  ( .A(\ctlif/N91 ), .B(\ctlif/N114 ), .Z(\ctlif/N115 ) );
  GTECH_OR2 \ctlif/C1640  ( .A(\ctlif/N88 ), .B(\ctlif/N113 ), .Z(\ctlif/N114 ) );
  GTECH_OR2 \ctlif/C1639  ( .A(\ctlif/N86 ), .B(\ctlif/N112 ), .Z(\ctlif/N113 ) );
  GTECH_OR2 \ctlif/C1638  ( .A(\ctlif/N83 ), .B(\ctlif/N111 ), .Z(\ctlif/N112 ) );
  GTECH_OR2 \ctlif/C1637  ( .A(\ctlif/N81 ), .B(\ctlif/N110 ), .Z(\ctlif/N111 ) );
  GTECH_OR2 \ctlif/C1636  ( .A(\ctlif/N79 ), .B(\ctlif/N109 ), .Z(\ctlif/N110 ) );
  GTECH_OR2 \ctlif/C1635  ( .A(\ctlif/N77 ), .B(\ctlif/N108 ), .Z(\ctlif/N109 ) );
  GTECH_OR2 \ctlif/C1634  ( .A(\ctlif/N74 ), .B(\ctlif/N107 ), .Z(\ctlif/N108 ) );
  GTECH_OR2 \ctlif/C1633  ( .A(\ctlif/N72 ), .B(\ctlif/N70 ), .Z(\ctlif/N107 )
         );
  GTECH_NOT \ctlif/I_21  ( .A(\ctlif/N105 ), .Z(\ctlif/N106 ) );
  GTECH_NOT \ctlif/I_20  ( .A(csr_a[2]), .Z(\ctlif/N102 ) );
  GTECH_NOT \ctlif/I_19  ( .A(csr_a[3]), .Z(\ctlif/N101 ) );
  GTECH_NOT \ctlif/I_18  ( .A(\ctlif/N99 ), .Z(\ctlif/N100 ) );
  GTECH_NOT \ctlif/I_17  ( .A(csr_a[0]), .Z(\ctlif/N96 ) );
  GTECH_NOT \ctlif/I_16  ( .A(csr_a[1]), .Z(\ctlif/N95 ) );
  GTECH_NOT \ctlif/I_15  ( .A(\ctlif/N93 ), .Z(\ctlif/N94 ) );
  GTECH_NOT \ctlif/I_14  ( .A(\ctlif/N90 ), .Z(\ctlif/N91 ) );
  GTECH_NOT \ctlif/I_13  ( .A(\ctlif/N87 ), .Z(\ctlif/N88 ) );
  GTECH_NOT \ctlif/I_12  ( .A(\ctlif/N85 ), .Z(\ctlif/N86 ) );
  GTECH_NOT \ctlif/I_11  ( .A(\ctlif/N82 ), .Z(\ctlif/N83 ) );
  GTECH_NOT \ctlif/I_10  ( .A(\ctlif/N80 ), .Z(\ctlif/N81 ) );
  GTECH_NOT \ctlif/I_9  ( .A(\ctlif/N78 ), .Z(\ctlif/N79 ) );
  GTECH_NOT \ctlif/I_8  ( .A(\ctlif/N76 ), .Z(\ctlif/N77 ) );
  GTECH_NOT \ctlif/I_7  ( .A(\ctlif/N73 ), .Z(\ctlif/N74 ) );
  GTECH_NOT \ctlif/I_6  ( .A(\ctlif/N71 ), .Z(\ctlif/N72 ) );
  GTECH_NOT \ctlif/I_5  ( .A(csr_we), .Z(\ctlif/N55 ) );
  GTECH_NOT \ctlif/I_4  ( .A(sys_rst), .Z(\ctlif/N54 ) );
  GTECH_AND2 \ctlif/C1594  ( .A(baseaddress_ack), .B(\ctlif/N52 ), .Z(
        \ctlif/N53 ) );
  GTECH_NOT \ctlif/I_3  ( .A(sys_rst), .Z(\ctlif/N52 ) );
  GTECH_NOT \ctlif/I_2  ( .A(\ctlif/sda_o ), .Z(\ctlif/N272 ) );
  GTECH_AND2 \ctlif/C1587  ( .A(\ctlif/sda_oe ), .B(\ctlif/N272 ), .Z(
        \ctlif/N24 ) );
  SELECT_OP \ctlif/C1584  ( .DATA1(1'b1), .DATA2(\ctlif/N146 ), .CONTROL1(
        \ctlif/N1 ), .CONTROL2(\ctlif/N23 ), .Z(\ctlif/N259 ) );
  SELECT_OP \ctlif/C1583  ( .DATA1(1'b1), .DATA2(\ctlif/N157 ), .CONTROL1(
        \ctlif/N1 ), .CONTROL2(\ctlif/N23 ), .Z(\ctlif/N258 ) );
  SELECT_OP \ctlif/C1582  ( .DATA1({1'b1, 1'b1}), .DATA2({csr_di[14], 
        csr_di[11]}), .CONTROL1(\ctlif/N1 ), .CONTROL2(\ctlif/N23 ), .Z({
        \ctlif/N257 , \ctlif/N256 }) );
  SELECT_OP \ctlif/C1581  ( .DATA1(1'b1), .DATA2(\ctlif/N156 ), .CONTROL1(
        \ctlif/N1 ), .CONTROL2(\ctlif/N23 ), .Z(\ctlif/N255 ) );
  SELECT_OP \ctlif/C1580  ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .DATA2(csr_di[25:11]), .CONTROL1(\ctlif/N1 ), .CONTROL2(\ctlif/N23 ), .Z({\ctlif/N254 , 
        \ctlif/N253 , \ctlif/N252 , \ctlif/N251 , \ctlif/N250 , \ctlif/N249 , 
        \ctlif/N248 , \ctlif/N247 , \ctlif/N246 , \ctlif/N245 , \ctlif/N244 , 
        \ctlif/N243 , \ctlif/N242 , \ctlif/N241 , \ctlif/N240 }) );
  SELECT_OP \ctlif/C1579  ( .DATA1(1'b1), .DATA2(\ctlif/N155 ), .CONTROL1(
        \ctlif/N1 ), .CONTROL2(\ctlif/N23 ), .Z(\ctlif/N239 ) );
  SELECT_OP \ctlif/C1578  ( .DATA1(1'b1), .DATA2(\ctlif/N154 ), .CONTROL1(
        \ctlif/N1 ), .CONTROL2(\ctlif/N23 ), .Z(\ctlif/N238 ) );
  SELECT_OP \ctlif/C1577  ( .DATA1(1'b1), .DATA2(\ctlif/N153 ), .CONTROL1(
        \ctlif/N1 ), .CONTROL2(\ctlif/N23 ), .Z(\ctlif/N237 ) );
  SELECT_OP \ctlif/C1576  ( .DATA1(1'b1), .DATA2(\ctlif/N152 ), .CONTROL1(
        \ctlif/N1 ), .CONTROL2(\ctlif/N23 ), .Z(\ctlif/N236 ) );
  SELECT_OP \ctlif/C1575  ( .DATA1(1'b0), .DATA2(csr_di[9]), .CONTROL1(
        \ctlif/N1 ), .CONTROL2(\ctlif/N23 ), .Z(\ctlif/N235 ) );
  SELECT_OP \ctlif/C1574  ( .DATA1(1'b1), .DATA2(\ctlif/N151 ), .CONTROL1(
        \ctlif/N1 ), .CONTROL2(\ctlif/N23 ), .Z(\ctlif/N234 ) );
  SELECT_OP \ctlif/C1573  ( .DATA1({1'b1, 1'b0, 1'b1, 1'b1, 1'b1}), .DATA2({
        csr_di[8:7], csr_di[3:1]}), .CONTROL1(\ctlif/N1 ), .CONTROL2(
        \ctlif/N23 ), .Z({\ctlif/N233 , \ctlif/N232 , \ctlif/N231 , 
        \ctlif/N230 , \ctlif/N229 }) );
  SELECT_OP \ctlif/C1572  ( .DATA1(1'b1), .DATA2(\ctlif/N150 ), .CONTROL1(
        \ctlif/N1 ), .CONTROL2(\ctlif/N23 ), .Z(\ctlif/N228 ) );
  SELECT_OP \ctlif/C1571  ( .DATA1({1'b1, 1'b1}), .DATA2(csr_di[6:5]), 
        .CONTROL1(\ctlif/N1 ), .CONTROL2(\ctlif/N23 ), .Z({\ctlif/N227 , 
        \ctlif/N226 }) );
  SELECT_OP \ctlif/C1570  ( .DATA1(1'b1), .DATA2(\ctlif/N149 ), .CONTROL1(
        \ctlif/N1 ), .CONTROL2(\ctlif/N23 ), .Z(\ctlif/N225 ) );
  SELECT_OP \ctlif/C1569  ( .DATA1(1'b1), .DATA2(csr_di[4]), .CONTROL1(
        \ctlif/N1 ), .CONTROL2(\ctlif/N23 ), .Z(\ctlif/N224 ) );
  SELECT_OP \ctlif/C1568  ( .DATA1(1'b1), .DATA2(\ctlif/N148 ), .CONTROL1(
        \ctlif/N1 ), .CONTROL2(\ctlif/N23 ), .Z(\ctlif/N223 ) );
  SELECT_OP \ctlif/C1567  ( .DATA1({1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .DATA2(csr_di[10:0]), .CONTROL1(\ctlif/N1 ), 
        .CONTROL2(\ctlif/N23 ), .Z({\ctlif/N222 , \ctlif/N221 , \ctlif/N220 , 
        \ctlif/N219 , \ctlif/N218 , \ctlif/N217 , \ctlif/N216 , \ctlif/N215 , 
        \ctlif/N214 , \ctlif/N213 , \ctlif/N212 }) );
  SELECT_OP \ctlif/C1566  ( .DATA1(1'b1), .DATA2(\ctlif/N147 ), .CONTROL1(
        \ctlif/N1 ), .CONTROL2(\ctlif/N23 ), .Z(\ctlif/N211 ) );
  SELECT_OP \ctlif/C1565  ( .DATA1(1'b1), .DATA2(csr_di[0]), .CONTROL1(
        \ctlif/N1 ), .CONTROL2(\ctlif/N23 ), .Z(\ctlif/N210 ) );
  GTECH_BUF \ctlif/B_22  ( .A(\ctlif/N54 ), .Z(\ctlif/N23 ) );
  SELECT_OP \ctlif/C1564  ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .DATA2({\ctlif/N183 , 
        \ctlif/N182 , \ctlif/N181 , \ctlif/N180 , \ctlif/N179 , \ctlif/N178 , 
        \ctlif/N177 , \ctlif/N176 , \ctlif/N175 , \ctlif/N174 , \ctlif/N173 , 
        \ctlif/N172 , \ctlif/N171 , \ctlif/N170 , \ctlif/N169 , \ctlif/N168 , 
        \ctlif/N167 , \ctlif/N166 , \ctlif/N165 , \ctlif/N164 , \ctlif/N163 , 
        \ctlif/N162 , \ctlif/N161 , \ctlif/N160 , \ctlif/N159 , \ctlif/N158 }), 
        .CONTROL1(\ctlif/N1 ), .CONTROL2(\ctlif/N23 ), .Z({\ctlif/N209 , 
        \ctlif/N208 , \ctlif/N207 , \ctlif/N206 , \ctlif/N205 , \ctlif/N204 , 
        \ctlif/N203 , \ctlif/N202 , \ctlif/N201 , \ctlif/N200 , \ctlif/N199 , 
        \ctlif/N198 , \ctlif/N197 , \ctlif/N196 , \ctlif/N195 , \ctlif/N194 , 
        \ctlif/N193 , \ctlif/N192 , \ctlif/N191 , \ctlif/N190 , \ctlif/N189 , 
        \ctlif/N188 , \ctlif/N187 , \ctlif/N186 , \ctlif/N185 , \ctlif/N184 })
         );
  SELECT_OP \ctlif/C1563  ( .DATA1({\ctlif/N145 , \ctlif/N144 , \ctlif/N143 , 
        \ctlif/N142 , \ctlif/N141 , \ctlif/N140 , \ctlif/N139 , \ctlif/N138 , 
        \ctlif/N137 , \ctlif/N136 , \ctlif/N135 , \ctlif/N134 , \ctlif/N133 , 
        \ctlif/N132 , \ctlif/N131 , \ctlif/N130 , \ctlif/N129 , \ctlif/N128 , 
        \ctlif/N127 , \ctlif/N126 , \ctlif/N125 , \ctlif/N124 , \ctlif/N123 , 
        \ctlif/N122 , \ctlif/N121 , \ctlif/N120 }), .DATA2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .CONTROL1(\ctlif/N21 ), .CONTROL2(\ctlif/N22 ), .Z({\ctlif/N183 , 
        \ctlif/N182 , \ctlif/N181 , \ctlif/N180 , \ctlif/N179 , \ctlif/N178 , 
        \ctlif/N177 , \ctlif/N176 , \ctlif/N175 , \ctlif/N174 , \ctlif/N173 , 
        \ctlif/N172 , \ctlif/N171 , \ctlif/N170 , \ctlif/N169 , \ctlif/N168 , 
        \ctlif/N167 , \ctlif/N166 , \ctlif/N165 , \ctlif/N164 , \ctlif/N163 , 
        \ctlif/N162 , \ctlif/N161 , \ctlif/N160 , \ctlif/N159 , \ctlif/N158 })
         );
  SELECT_OP \ctlif/C1562  ( .DATA1(\ctlif/N67 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N21 ), .CONTROL2(\ctlif/N22 ), .Z(\ctlif/N157 ) );
  SELECT_OP \ctlif/C1561  ( .DATA1(\ctlif/N66 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N21 ), .CONTROL2(\ctlif/N22 ), .Z(\ctlif/N156 ) );
  SELECT_OP \ctlif/C1560  ( .DATA1(\ctlif/N65 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N21 ), .CONTROL2(\ctlif/N22 ), .Z(\ctlif/N155 ) );
  SELECT_OP \ctlif/C1559  ( .DATA1(\ctlif/N64 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N21 ), .CONTROL2(\ctlif/N22 ), .Z(\ctlif/N154 ) );
  SELECT_OP \ctlif/C1558  ( .DATA1(\ctlif/N63 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N21 ), .CONTROL2(\ctlif/N22 ), .Z(\ctlif/N153 ) );
  SELECT_OP \ctlif/C1557  ( .DATA1(\ctlif/N62 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N21 ), .CONTROL2(\ctlif/N22 ), .Z(\ctlif/N152 ) );
  SELECT_OP \ctlif/C1556  ( .DATA1(\ctlif/N61 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N21 ), .CONTROL2(\ctlif/N22 ), .Z(\ctlif/N151 ) );
  SELECT_OP \ctlif/C1555  ( .DATA1(\ctlif/N60 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N21 ), .CONTROL2(\ctlif/N22 ), .Z(\ctlif/N150 ) );
  SELECT_OP \ctlif/C1554  ( .DATA1(\ctlif/N59 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N21 ), .CONTROL2(\ctlif/N22 ), .Z(\ctlif/N149 ) );
  SELECT_OP \ctlif/C1553  ( .DATA1(\ctlif/N58 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N21 ), .CONTROL2(\ctlif/N22 ), .Z(\ctlif/N148 ) );
  SELECT_OP \ctlif/C1552  ( .DATA1(\ctlif/N57 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N21 ), .CONTROL2(\ctlif/N22 ), .Z(\ctlif/N147 ) );
  GTECH_BUF \ctlif/B_21  ( .A(\ctlif/N262 ), .Z(\ctlif/N22 ) );
  GTECH_BUF \ctlif/B_20  ( .A(\ctlif/N263 ), .Z(\ctlif/N21 ) );
  SELECT_OP \ctlif/C1551  ( .DATA1(\ctlif/N56 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N21 ), .CONTROL2(\ctlif/N22 ), .Z(\ctlif/N146 ) );
  GTECH_BUF \ctlif/B_19  ( .A(\ctlif/N271 ), .Z(\ctlif/N20 ) );
  SELECT_OP \ctlif/C1550  ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .DATA2(baseaddress[25:18]), .DATA3(
        \ctlif/baseaddress_act [25:18]), .CONTROL1(\ctlif/N20 ), .CONTROL2(
        \ctlif/N13 ), .CONTROL3(\ctlif/N14 ), .Z({\ctlif/N145 , \ctlif/N144 , 
        \ctlif/N143 , \ctlif/N142 , \ctlif/N141 , \ctlif/N140 , \ctlif/N139 , 
        \ctlif/N138 }) );
  GTECH_BUF \ctlif/B_18  ( .A(\ctlif/N268 ), .Z(\ctlif/N19 ) );
  SELECT_OP \ctlif/C1549  ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(baseaddress[17:11]), .DATA3(\ctlif/baseaddress_act [17:11]), 
        .DATA4(nbursts[17:11]), .CONTROL1(\ctlif/N19 ), .CONTROL2(\ctlif/N13 ), 
        .CONTROL3(\ctlif/N14 ), .CONTROL4(\ctlif/N15 ), .Z({\ctlif/N137 , 
        \ctlif/N136 , \ctlif/N135 , \ctlif/N134 , \ctlif/N133 , \ctlif/N132 , 
        \ctlif/N131 }) );
  GTECH_BUF \ctlif/B_17  ( .A(\ctlif/N265 ), .Z(\ctlif/N18 ) );
  SELECT_OP \ctlif/C1548  ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(hres[10:4]), .DATA3(hsync_start[10:4]), .DATA4(hsync_end[10:4]), 
        .DATA5(hscan[10:4]), .DATA6(vres[10:4]), .DATA7(vsync_start[10:4]), 
        .DATA8(vsync_end[10:4]), .DATA9(vscan[10:4]), .DATA10(
        baseaddress[10:4]), .DATA11(\ctlif/baseaddress_act [10:4]), .DATA12(
        nbursts[10:4]), .CONTROL1(\ctlif/N18 ), .CONTROL2(\ctlif/N5 ), 
        .CONTROL3(\ctlif/N6 ), .CONTROL4(\ctlif/N7 ), .CONTROL5(\ctlif/N8 ), 
        .CONTROL6(\ctlif/N9 ), .CONTROL7(\ctlif/N10 ), .CONTROL8(\ctlif/N11 ), 
        .CONTROL9(\ctlif/N12 ), .CONTROL10(\ctlif/N13 ), .CONTROL11(
        \ctlif/N14 ), .CONTROL12(\ctlif/N15 ), .Z({\ctlif/N130 , \ctlif/N129 , 
        \ctlif/N128 , \ctlif/N127 , \ctlif/N126 , \ctlif/N125 , \ctlif/N124 })
         );
  GTECH_BUF \ctlif/B_16  ( .A(\ctlif/N264 ), .Z(\ctlif/N17 ) );
  SELECT_OP \ctlif/C1547  ( .DATA1({1'b0, 1'b0, 1'b0}), .DATA2(hres[3:1]), 
        .DATA3(hsync_start[3:1]), .DATA4(hsync_end[3:1]), .DATA5(hscan[3:1]), 
        .DATA6(vres[3:1]), .DATA7(vsync_start[3:1]), .DATA8(vsync_end[3:1]), 
        .DATA9(vscan[3:1]), .DATA10(baseaddress[3:1]), .DATA11(
        \ctlif/baseaddress_act [3:1]), .DATA12(nbursts[3:1]), .DATA13({vga_sdc, 
        \ctlif/sda_oe , \ctlif/sda_o }), .CONTROL1(\ctlif/N17 ), .CONTROL2(
        \ctlif/N5 ), .CONTROL3(\ctlif/N6 ), .CONTROL4(\ctlif/N7 ), .CONTROL5(
        \ctlif/N8 ), .CONTROL6(\ctlif/N9 ), .CONTROL7(\ctlif/N10 ), .CONTROL8(
        \ctlif/N11 ), .CONTROL9(\ctlif/N12 ), .CONTROL10(\ctlif/N13 ), 
        .CONTROL11(\ctlif/N14 ), .CONTROL12(\ctlif/N15 ), .CONTROL13(
        \ctlif/N16 ), .Z({\ctlif/N123 , \ctlif/N122 , \ctlif/N121 }) );
  GTECH_BUF \ctlif/B_15  ( .A(\ctlif/N106 ), .Z(\ctlif/N16 ) );
  GTECH_BUF \ctlif/B_14  ( .A(\ctlif/N100 ), .Z(\ctlif/N15 ) );
  GTECH_BUF \ctlif/B_13  ( .A(\ctlif/N94 ), .Z(\ctlif/N14 ) );
  GTECH_BUF \ctlif/B_12  ( .A(\ctlif/N91 ), .Z(\ctlif/N13 ) );
  GTECH_BUF \ctlif/B_11  ( .A(\ctlif/N88 ), .Z(\ctlif/N12 ) );
  GTECH_BUF \ctlif/B_10  ( .A(\ctlif/N86 ), .Z(\ctlif/N11 ) );
  GTECH_BUF \ctlif/B_9  ( .A(\ctlif/N83 ), .Z(\ctlif/N10 ) );
  GTECH_BUF \ctlif/B_8  ( .A(\ctlif/N81 ), .Z(\ctlif/N9 ) );
  GTECH_BUF \ctlif/B_7  ( .A(\ctlif/N79 ), .Z(\ctlif/N8 ) );
  GTECH_BUF \ctlif/B_6  ( .A(\ctlif/N77 ), .Z(\ctlif/N7 ) );
  GTECH_BUF \ctlif/B_5  ( .A(\ctlif/N74 ), .Z(\ctlif/N6 ) );
  GTECH_BUF \ctlif/B_4  ( .A(\ctlif/N72 ), .Z(\ctlif/N5 ) );
  GTECH_BUF \ctlif/B_3  ( .A(\ctlif/N70 ), .Z(\ctlif/N4 ) );
  SELECT_OP \ctlif/C1546  ( .DATA1(vga_rst), .DATA2(hres[0]), .DATA3(
        hsync_start[0]), .DATA4(hsync_end[0]), .DATA5(hscan[0]), .DATA6(
        vres[0]), .DATA7(vsync_start[0]), .DATA8(vsync_end[0]), .DATA9(
        vscan[0]), .DATA10(baseaddress[0]), .DATA11(\ctlif/baseaddress_act [0]), .DATA12(nbursts[0]), .DATA13(\ctlif/sda_2 ), .DATA14(1'b0), .CONTROL1(
        \ctlif/N4 ), .CONTROL2(\ctlif/N5 ), .CONTROL3(\ctlif/N6 ), .CONTROL4(
        \ctlif/N7 ), .CONTROL5(\ctlif/N8 ), .CONTROL6(\ctlif/N9 ), .CONTROL7(
        \ctlif/N10 ), .CONTROL8(\ctlif/N11 ), .CONTROL9(\ctlif/N12 ), 
        .CONTROL10(\ctlif/N13 ), .CONTROL11(\ctlif/N14 ), .CONTROL12(
        \ctlif/N15 ), .CONTROL13(\ctlif/N16 ), .CONTROL14(\ctlif/N119 ), .Z(
        \ctlif/N120 ) );
  SELECT_OP \ctlif/C1545  ( .DATA1(\ctlif/N100 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N2 ), .CONTROL2(\ctlif/N3 ), .Z(\ctlif/N67 ) );
  SELECT_OP \ctlif/C1544  ( .DATA1(\ctlif/N91 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N2 ), .CONTROL2(\ctlif/N3 ), .Z(\ctlif/N66 ) );
  SELECT_OP \ctlif/C1543  ( .DATA1(\ctlif/N88 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N2 ), .CONTROL2(\ctlif/N3 ), .Z(\ctlif/N65 ) );
  SELECT_OP \ctlif/C1542  ( .DATA1(\ctlif/N86 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N2 ), .CONTROL2(\ctlif/N3 ), .Z(\ctlif/N64 ) );
  SELECT_OP \ctlif/C1541  ( .DATA1(\ctlif/N83 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N2 ), .CONTROL2(\ctlif/N3 ), .Z(\ctlif/N63 ) );
  SELECT_OP \ctlif/C1540  ( .DATA1(\ctlif/N81 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N2 ), .CONTROL2(\ctlif/N3 ), .Z(\ctlif/N62 ) );
  SELECT_OP \ctlif/C1539  ( .DATA1(\ctlif/N79 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N2 ), .CONTROL2(\ctlif/N3 ), .Z(\ctlif/N61 ) );
  SELECT_OP \ctlif/C1538  ( .DATA1(\ctlif/N77 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N2 ), .CONTROL2(\ctlif/N3 ), .Z(\ctlif/N60 ) );
  SELECT_OP \ctlif/C1537  ( .DATA1(\ctlif/N74 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N2 ), .CONTROL2(\ctlif/N3 ), .Z(\ctlif/N59 ) );
  SELECT_OP \ctlif/C1536  ( .DATA1(\ctlif/N72 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N2 ), .CONTROL2(\ctlif/N3 ), .Z(\ctlif/N58 ) );
  SELECT_OP \ctlif/C1535  ( .DATA1(\ctlif/N70 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N2 ), .CONTROL2(\ctlif/N3 ), .Z(\ctlif/N57 ) );
  GTECH_BUF \ctlif/B_2  ( .A(\ctlif/N55 ), .Z(\ctlif/N3 ) );
  GTECH_BUF \ctlif/B_1  ( .A(csr_we), .Z(\ctlif/N2 ) );
  SELECT_OP \ctlif/C1534  ( .DATA1(\ctlif/N106 ), .DATA2(1'b0), .CONTROL1(
        \ctlif/N2 ), .CONTROL2(\ctlif/N3 ), .Z(\ctlif/N56 ) );
  GTECH_BUF \ctlif/B_0  ( .A(sys_rst), .Z(\ctlif/N1 ) );
  SELECT_OP \ctlif/C1533  ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .DATA2(baseaddress), 
        .CONTROL1(\ctlif/N1 ), .CONTROL2(\ctlif/N53 ), .Z({\ctlif/N51 , 
        \ctlif/N50 , \ctlif/N49 , \ctlif/N48 , \ctlif/N47 , \ctlif/N46 , 
        \ctlif/N45 , \ctlif/N44 , \ctlif/N43 , \ctlif/N42 , \ctlif/N41 , 
        \ctlif/N40 , \ctlif/N39 , \ctlif/N38 , \ctlif/N37 , \ctlif/N36 , 
        \ctlif/N35 , \ctlif/N34 , \ctlif/N33 , \ctlif/N32 , \ctlif/N31 , 
        \ctlif/N30 , \ctlif/N29 , \ctlif/N28 , \ctlif/N27 , \ctlif/N26 }) );
  GTECH_OR3 \ctlif/C1495  ( .A(\ctlif/N266 ), .B(\ctlif/N269 ), .C(
        \ctlif/N270 ), .Z(\ctlif/N271 ) );
  GTECH_OR2 \ctlif/C1494  ( .A(\ctlif/N106 ), .B(\ctlif/N119 ), .Z(
        \ctlif/N270 ) );
  GTECH_OR5 \ctlif/C1493  ( .A(\ctlif/N81 ), .B(\ctlif/N83 ), .C(\ctlif/N86 ), 
        .D(\ctlif/N88 ), .E(\ctlif/N100 ), .Z(\ctlif/N269 ) );
  GTECH_OR3 \ctlif/C1466  ( .A(\ctlif/N266 ), .B(\ctlif/N267 ), .C(
        \ctlif/N119 ), .Z(\ctlif/N268 ) );
  GTECH_OR5 \ctlif/C1465  ( .A(\ctlif/N81 ), .B(\ctlif/N83 ), .C(\ctlif/N86 ), 
        .D(\ctlif/N88 ), .E(\ctlif/N106 ), .Z(\ctlif/N267 ) );
  GTECH_OR5 \ctlif/C1464  ( .A(\ctlif/N70 ), .B(\ctlif/N72 ), .C(\ctlif/N74 ), 
        .D(\ctlif/N77 ), .E(\ctlif/N79 ), .Z(\ctlif/N266 ) );
  GTECH_OR3 \ctlif/C1450  ( .A(\ctlif/N70 ), .B(\ctlif/N106 ), .C(\ctlif/N119 ), .Z(\ctlif/N265 ) );
  GTECH_OR2 \ctlif/C1444  ( .A(\ctlif/N70 ), .B(\ctlif/N119 ), .Z(\ctlif/N264 ) );
  GTECH_OR2 \ctlif/C1332  ( .A(sys_rst), .B(\ctlif/N53 ), .Z(\ctlif/N25 ) );
  GTECH_NOT \ctlif/I_1  ( .A(\ctlif/N262 ), .Z(\ctlif/N263 ) );
  GTECH_OR2 \ctlif/C1330  ( .A(csr_a[10]), .B(\ctlif/N261 ), .Z(\ctlif/N262 )
         );
  GTECH_OR2 \ctlif/C1329  ( .A(csr_a[11]), .B(\ctlif/N260 ), .Z(\ctlif/N261 )
         );
  GTECH_OR2 \ctlif/C1328  ( .A(csr_a[12]), .B(csr_a[13]), .Z(\ctlif/N260 ) );
  \**SEQGEN**  \ctlif/sda_oe_reg  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N214 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(\ctlif/sda_oe ), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N259 ) );
  \**SEQGEN**  \ctlif/baseaddress_reg_0_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N212 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[0]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_1_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N213 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[1]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_2_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N214 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[2]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_3_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N215 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[3]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_4_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N216 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[4]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_5_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N217 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[5]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_6_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N218 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[6]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_7_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N232 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[7]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_8_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N220 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[8]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_9_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N235 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[9]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_10_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N222 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[10]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_11_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N240 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[11]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_12_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N241 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[12]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_13_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N242 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[13]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_14_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N243 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[14]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_15_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N244 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[15]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_16_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N245 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[16]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_17_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N246 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[17]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_18_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N247 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[18]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_19_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N248 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[19]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_20_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N249 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[20]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_21_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N250 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[21]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_22_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N251 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[22]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_23_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N252 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[23]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_24_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N253 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[24]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/baseaddress_reg_25_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N254 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(baseaddress[25]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N255 )
         );
  \**SEQGEN**  \ctlif/vres_reg_0_  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N212 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(vres[0]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N236 ) );
  \**SEQGEN**  \ctlif/vres_reg_1_  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N213 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(vres[1]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N236 ) );
  \**SEQGEN**  \ctlif/vres_reg_2_  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N214 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(vres[2]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N236 ) );
  \**SEQGEN**  \ctlif/vres_reg_3_  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N215 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(vres[3]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N236 ) );
  \**SEQGEN**  \ctlif/vres_reg_4_  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N216 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(vres[4]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N236 ) );
  \**SEQGEN**  \ctlif/vres_reg_5_  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N226 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(vres[5]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N236 ) );
  \**SEQGEN**  \ctlif/vres_reg_6_  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N227 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(vres[6]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N236 ) );
  \**SEQGEN**  \ctlif/vres_reg_7_  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N219 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(vres[7]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N236 ) );
  \**SEQGEN**  \ctlif/vres_reg_8_  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N233 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(vres[8]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N236 ) );
  \**SEQGEN**  \ctlif/vres_reg_9_  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N235 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(vres[9]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N236 ) );
  \**SEQGEN**  \ctlif/vres_reg_10_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N222 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vres[10]), .QN(), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N236 ) );
  \**SEQGEN**  \ctlif/nbursts_reg_0_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N212 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(nbursts[0]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N258 )
         );
  \**SEQGEN**  \ctlif/nbursts_reg_1_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N213 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(nbursts[1]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N258 )
         );
  \**SEQGEN**  \ctlif/nbursts_reg_2_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N214 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(nbursts[2]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N258 )
         );
  \**SEQGEN**  \ctlif/nbursts_reg_3_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N215 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(nbursts[3]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N258 )
         );
  \**SEQGEN**  \ctlif/nbursts_reg_4_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N216 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(nbursts[4]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N258 )
         );
  \**SEQGEN**  \ctlif/nbursts_reg_5_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N217 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(nbursts[5]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N258 )
         );
  \**SEQGEN**  \ctlif/nbursts_reg_6_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N218 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(nbursts[6]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N258 )
         );
  \**SEQGEN**  \ctlif/nbursts_reg_7_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N232 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(nbursts[7]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N258 )
         );
  \**SEQGEN**  \ctlif/nbursts_reg_8_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N233 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(nbursts[8]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N258 )
         );
  \**SEQGEN**  \ctlif/nbursts_reg_9_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N221 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(nbursts[9]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N258 )
         );
  \**SEQGEN**  \ctlif/nbursts_reg_10_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N222 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(nbursts[10]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N258 )
         );
  \**SEQGEN**  \ctlif/nbursts_reg_11_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N256 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(nbursts[11]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N258 )
         );
  \**SEQGEN**  \ctlif/nbursts_reg_12_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N241 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(nbursts[12]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N258 )
         );
  \**SEQGEN**  \ctlif/nbursts_reg_13_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N242 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(nbursts[13]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N258 )
         );
  \**SEQGEN**  \ctlif/nbursts_reg_14_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N257 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(nbursts[14]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N258 )
         );
  \**SEQGEN**  \ctlif/nbursts_reg_15_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N244 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(nbursts[15]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N258 )
         );
  \**SEQGEN**  \ctlif/nbursts_reg_16_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N245 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(nbursts[16]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N258 )
         );
  \**SEQGEN**  \ctlif/nbursts_reg_17_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N246 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(nbursts[17]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N258 )
         );
  \**SEQGEN**  \ctlif/vga_rst_reg  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N210 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(vga_rst), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N211 ) );
  \**SEQGEN**  \ctlif/csr_do_reg_0_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N184 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[0]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_1_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N185 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[1]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_2_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N186 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[2]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_3_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N187 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[3]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_4_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N188 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[4]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_5_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N189 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[5]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_6_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N190 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[6]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_7_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N191 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[7]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_8_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N192 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[8]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_9_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N193 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[9]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_10_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N194 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[10]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_11_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N195 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[11]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_12_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N196 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[12]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_13_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N197 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[13]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_14_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N198 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[14]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_15_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N199 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[15]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_16_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N200 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[16]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_17_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N201 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[17]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_18_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N202 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[18]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_19_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N203 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[19]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_20_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N204 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[20]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_21_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N205 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[21]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_22_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N206 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[22]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_23_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N207 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[23]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_24_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N208 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[24]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_25_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N209 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(csr_do[25]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_26_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(csr_do[26]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_27_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(csr_do[27]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_28_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(csr_do[28]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_29_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(csr_do[29]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_30_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(csr_do[30]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/csr_do_reg_31_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(csr_do[31]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/hres_reg_0_  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N212 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(hres[0]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N223 ) );
  \**SEQGEN**  \ctlif/hres_reg_1_  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N213 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(hres[1]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N223 ) );
  \**SEQGEN**  \ctlif/hres_reg_2_  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N214 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(hres[2]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N223 ) );
  \**SEQGEN**  \ctlif/hres_reg_3_  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N215 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(hres[3]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N223 ) );
  \**SEQGEN**  \ctlif/hres_reg_4_  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N216 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(hres[4]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N223 ) );
  \**SEQGEN**  \ctlif/hres_reg_5_  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N217 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(hres[5]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N223 ) );
  \**SEQGEN**  \ctlif/hres_reg_6_  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N218 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(hres[6]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N223 ) );
  \**SEQGEN**  \ctlif/hres_reg_7_  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N219 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(hres[7]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N223 ) );
  \**SEQGEN**  \ctlif/hres_reg_8_  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N220 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(hres[8]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N223 ) );
  \**SEQGEN**  \ctlif/hres_reg_9_  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N221 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(hres[9]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N223 ) );
  \**SEQGEN**  \ctlif/hres_reg_10_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N222 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hres[10]), .QN(), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N223 ) );
  \**SEQGEN**  \ctlif/sda_o_reg  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N213 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(\ctlif/sda_o ), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N259 ) );
  \**SEQGEN**  \ctlif/vga_sdc_reg  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/N215 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(vga_sdc), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\ctlif/N259 ) );
  \**SEQGEN**  \ctlif/hsync_end_reg_0_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N212 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hsync_end[0]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N228 )
         );
  \**SEQGEN**  \ctlif/hsync_end_reg_1_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N213 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hsync_end[1]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N228 )
         );
  \**SEQGEN**  \ctlif/hsync_end_reg_2_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N214 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hsync_end[2]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N228 )
         );
  \**SEQGEN**  \ctlif/hsync_end_reg_3_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N215 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hsync_end[3]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N228 )
         );
  \**SEQGEN**  \ctlif/hsync_end_reg_4_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N224 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hsync_end[4]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N228 )
         );
  \**SEQGEN**  \ctlif/hsync_end_reg_5_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N226 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hsync_end[5]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N228 )
         );
  \**SEQGEN**  \ctlif/hsync_end_reg_6_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N227 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hsync_end[6]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N228 )
         );
  \**SEQGEN**  \ctlif/hsync_end_reg_7_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N219 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hsync_end[7]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N228 )
         );
  \**SEQGEN**  \ctlif/hsync_end_reg_8_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N220 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hsync_end[8]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N228 )
         );
  \**SEQGEN**  \ctlif/hsync_end_reg_9_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N221 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hsync_end[9]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N228 )
         );
  \**SEQGEN**  \ctlif/hsync_end_reg_10_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N222 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hsync_end[10]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N228 )
         );
  \**SEQGEN**  \ctlif/hsync_start_reg_0_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N212 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hsync_start[0]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N225 )
         );
  \**SEQGEN**  \ctlif/hsync_start_reg_1_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N213 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hsync_start[1]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N225 )
         );
  \**SEQGEN**  \ctlif/hsync_start_reg_2_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N214 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hsync_start[2]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N225 )
         );
  \**SEQGEN**  \ctlif/hsync_start_reg_3_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N215 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hsync_start[3]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N225 )
         );
  \**SEQGEN**  \ctlif/hsync_start_reg_4_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N224 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hsync_start[4]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N225 )
         );
  \**SEQGEN**  \ctlif/hsync_start_reg_5_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N217 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hsync_start[5]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N225 )
         );
  \**SEQGEN**  \ctlif/hsync_start_reg_6_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N218 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hsync_start[6]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N225 )
         );
  \**SEQGEN**  \ctlif/hsync_start_reg_7_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N219 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hsync_start[7]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N225 )
         );
  \**SEQGEN**  \ctlif/hsync_start_reg_8_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N220 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hsync_start[8]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N225 )
         );
  \**SEQGEN**  \ctlif/hsync_start_reg_9_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N221 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hsync_start[9]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N225 )
         );
  \**SEQGEN**  \ctlif/hsync_start_reg_10_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N222 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hsync_start[10]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N225 )
         );
  \**SEQGEN**  \ctlif/hscan_reg_0_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N210 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hscan[0]), .QN(), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N234 ) );
  \**SEQGEN**  \ctlif/hscan_reg_1_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N229 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hscan[1]), .QN(), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N234 ) );
  \**SEQGEN**  \ctlif/hscan_reg_2_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N230 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hscan[2]), .QN(), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N234 ) );
  \**SEQGEN**  \ctlif/hscan_reg_3_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N231 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hscan[3]), .QN(), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N234 ) );
  \**SEQGEN**  \ctlif/hscan_reg_4_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N224 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hscan[4]), .QN(), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N234 ) );
  \**SEQGEN**  \ctlif/hscan_reg_5_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N217 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hscan[5]), .QN(), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N234 ) );
  \**SEQGEN**  \ctlif/hscan_reg_6_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N218 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hscan[6]), .QN(), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N234 ) );
  \**SEQGEN**  \ctlif/hscan_reg_7_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N232 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hscan[7]), .QN(), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N234 ) );
  \**SEQGEN**  \ctlif/hscan_reg_8_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N233 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hscan[8]), .QN(), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N234 ) );
  \**SEQGEN**  \ctlif/hscan_reg_9_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N221 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hscan[9]), .QN(), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N234 ) );
  \**SEQGEN**  \ctlif/hscan_reg_10_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N222 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(hscan[10]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N234 )
         );
  \**SEQGEN**  \ctlif/vsync_start_reg_0_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N210 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vsync_start[0]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N237 )
         );
  \**SEQGEN**  \ctlif/vsync_start_reg_1_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N229 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vsync_start[1]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N237 )
         );
  \**SEQGEN**  \ctlif/vsync_start_reg_2_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N214 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vsync_start[2]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N237 )
         );
  \**SEQGEN**  \ctlif/vsync_start_reg_3_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N231 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vsync_start[3]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N237 )
         );
  \**SEQGEN**  \ctlif/vsync_start_reg_4_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N216 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vsync_start[4]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N237 )
         );
  \**SEQGEN**  \ctlif/vsync_start_reg_5_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N226 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vsync_start[5]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N237 )
         );
  \**SEQGEN**  \ctlif/vsync_start_reg_6_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N227 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vsync_start[6]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N237 )
         );
  \**SEQGEN**  \ctlif/vsync_start_reg_7_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N219 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vsync_start[7]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N237 )
         );
  \**SEQGEN**  \ctlif/vsync_start_reg_8_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N233 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vsync_start[8]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N237 )
         );
  \**SEQGEN**  \ctlif/vsync_start_reg_9_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N235 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vsync_start[9]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N237 )
         );
  \**SEQGEN**  \ctlif/vsync_start_reg_10_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N222 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vsync_start[10]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N237 )
         );
  \**SEQGEN**  \ctlif/vsync_end_reg_0_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N210 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vsync_end[0]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N238 )
         );
  \**SEQGEN**  \ctlif/vsync_end_reg_1_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N213 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vsync_end[1]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N238 )
         );
  \**SEQGEN**  \ctlif/vsync_end_reg_2_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N230 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vsync_end[2]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N238 )
         );
  \**SEQGEN**  \ctlif/vsync_end_reg_3_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N231 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vsync_end[3]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N238 )
         );
  \**SEQGEN**  \ctlif/vsync_end_reg_4_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N216 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vsync_end[4]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N238 )
         );
  \**SEQGEN**  \ctlif/vsync_end_reg_5_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N226 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vsync_end[5]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N238 )
         );
  \**SEQGEN**  \ctlif/vsync_end_reg_6_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N227 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vsync_end[6]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N238 )
         );
  \**SEQGEN**  \ctlif/vsync_end_reg_7_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N219 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vsync_end[7]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N238 )
         );
  \**SEQGEN**  \ctlif/vsync_end_reg_8_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N233 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vsync_end[8]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N238 )
         );
  \**SEQGEN**  \ctlif/vsync_end_reg_9_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N235 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vsync_end[9]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N238 )
         );
  \**SEQGEN**  \ctlif/vsync_end_reg_10_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N222 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vsync_end[10]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N238 )
         );
  \**SEQGEN**  \ctlif/vscan_reg_0_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N210 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vscan[0]), .QN(), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N239 ) );
  \**SEQGEN**  \ctlif/vscan_reg_1_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N229 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vscan[1]), .QN(), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N239 ) );
  \**SEQGEN**  \ctlif/vscan_reg_2_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N214 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vscan[2]), .QN(), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N239 ) );
  \**SEQGEN**  \ctlif/vscan_reg_3_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N231 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vscan[3]), .QN(), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N239 ) );
  \**SEQGEN**  \ctlif/vscan_reg_4_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N216 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vscan[4]), .QN(), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N239 ) );
  \**SEQGEN**  \ctlif/vscan_reg_5_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N217 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vscan[5]), .QN(), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N239 ) );
  \**SEQGEN**  \ctlif/vscan_reg_6_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N218 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vscan[6]), .QN(), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N239 ) );
  \**SEQGEN**  \ctlif/vscan_reg_7_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N232 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vscan[7]), .QN(), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N239 ) );
  \**SEQGEN**  \ctlif/vscan_reg_8_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N220 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vscan[8]), .QN(), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N239 ) );
  \**SEQGEN**  \ctlif/vscan_reg_9_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N221 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vscan[9]), .QN(), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N239 ) );
  \**SEQGEN**  \ctlif/vscan_reg_10_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N222 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(vscan[10]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(\ctlif/N239 )
         );
  GTECH_OR2 \ctlif/C569  ( .A(\ctlif/N103 ), .B(\ctlif/N104 ), .Z(\ctlif/N105 ) );
  GTECH_OR2 \ctlif/C568  ( .A(csr_a[1]), .B(csr_a[0]), .Z(\ctlif/N104 ) );
  GTECH_OR2 \ctlif/C567  ( .A(\ctlif/N101 ), .B(\ctlif/N102 ), .Z(\ctlif/N103 ) );
  GTECH_OR2 \ctlif/C563  ( .A(\ctlif/N97 ), .B(\ctlif/N98 ), .Z(\ctlif/N99 )
         );
  GTECH_OR2 \ctlif/C562  ( .A(\ctlif/N95 ), .B(\ctlif/N96 ), .Z(\ctlif/N98 )
         );
  GTECH_OR2 \ctlif/C561  ( .A(\ctlif/N101 ), .B(csr_a[2]), .Z(\ctlif/N97 ) );
  GTECH_OR2 \ctlif/C556  ( .A(\ctlif/N97 ), .B(\ctlif/N92 ), .Z(\ctlif/N93 )
         );
  GTECH_OR2 \ctlif/C555  ( .A(\ctlif/N95 ), .B(csr_a[0]), .Z(\ctlif/N92 ) );
  GTECH_OR2 \ctlif/C550  ( .A(\ctlif/N97 ), .B(\ctlif/N89 ), .Z(\ctlif/N90 )
         );
  GTECH_OR2 \ctlif/C549  ( .A(csr_a[1]), .B(\ctlif/N96 ), .Z(\ctlif/N89 ) );
  GTECH_OR2 \ctlif/C544  ( .A(\ctlif/N97 ), .B(\ctlif/N104 ), .Z(\ctlif/N87 )
         );
  GTECH_OR2 \ctlif/C539  ( .A(\ctlif/N84 ), .B(\ctlif/N98 ), .Z(\ctlif/N85 )
         );
  GTECH_OR2 \ctlif/C537  ( .A(csr_a[3]), .B(\ctlif/N102 ), .Z(\ctlif/N84 ) );
  GTECH_OR2 \ctlif/C532  ( .A(\ctlif/N84 ), .B(\ctlif/N92 ), .Z(\ctlif/N82 )
         );
  GTECH_OR2 \ctlif/C526  ( .A(\ctlif/N84 ), .B(\ctlif/N89 ), .Z(\ctlif/N80 )
         );
  GTECH_OR2 \ctlif/C520  ( .A(\ctlif/N84 ), .B(\ctlif/N104 ), .Z(\ctlif/N78 )
         );
  GTECH_OR2 \ctlif/C515  ( .A(\ctlif/N75 ), .B(\ctlif/N98 ), .Z(\ctlif/N76 )
         );
  GTECH_OR2 \ctlif/C513  ( .A(csr_a[3]), .B(csr_a[2]), .Z(\ctlif/N75 ) );
  GTECH_OR2 \ctlif/C509  ( .A(\ctlif/N75 ), .B(\ctlif/N92 ), .Z(\ctlif/N73 )
         );
  GTECH_OR2 \ctlif/C504  ( .A(\ctlif/N75 ), .B(\ctlif/N89 ), .Z(\ctlif/N71 )
         );
  GTECH_AND2 \ctlif/C500  ( .A(\ctlif/N68 ), .B(\ctlif/N69 ), .Z(\ctlif/N70 )
         );
  GTECH_AND2 \ctlif/C499  ( .A(\ctlif/N95 ), .B(\ctlif/N96 ), .Z(\ctlif/N69 )
         );
  GTECH_AND2 \ctlif/C498  ( .A(\ctlif/N101 ), .B(\ctlif/N102 ), .Z(\ctlif/N68 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_0_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N26 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [0]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_1_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N27 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [1]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_2_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N28 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [2]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_3_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N29 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [3]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_4_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N30 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [4]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_5_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N31 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [5]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_6_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N32 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [6]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_7_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N33 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [7]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_8_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N34 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [8]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_9_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N35 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [9]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_10_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N36 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [10]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_11_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N37 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [11]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_12_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N38 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [12]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_13_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N39 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [13]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_14_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N40 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [14]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_15_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N41 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [15]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_16_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N42 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [16]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_17_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N43 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [17]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_18_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N44 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [18]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_19_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N45 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [19]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_20_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N46 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [20]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_21_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N47 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [21]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_22_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N48 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [22]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_23_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N49 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [23]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_24_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N50 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [24]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  \**SEQGEN**  \ctlif/baseaddress_act_reg_25_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\ctlif/N51 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\ctlif/baseaddress_act [25]), .QN(), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \ctlif/N25 ) );
  GTECH_NOT \ctlif/I_0  ( .A(\ctlif/N24 ), .Z(\ctlif/N0 ) );
  \**TSGEN**  \ctlif/vga_sda_tri  ( .\function (1'b0), .three_state(\ctlif/N0 ), .\output (vga_sda) );
  \**SEQGEN**  \ctlif/sda_2_reg  ( .clear(1'b0), .preset(1'b0), .next_state(
        \ctlif/sda_1 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(\ctlif/sda_2 ), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \ctlif/sda_1_reg  ( .clear(1'b0), .preset(1'b0), .next_state(
        vga_sda), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \ctlif/sda_1 ), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  GTECH_OR2 \pixelfeed/C705  ( .A(\pixelfeed/N40 ), .B(\pixelfeed/N245 ), .Z()
         );
  GTECH_AND2 \pixelfeed/C704  ( .A(\pixelfeed/N39 ), .B(\pixelfeed/N62 ), .Z(
        \pixelfeed/N246 ) );
  GTECH_OR2 \pixelfeed/C703  ( .A(\pixelfeed/N38 ), .B(\pixelfeed/N36 ), .Z(
        \pixelfeed/N245 ) );
  GTECH_NOT \pixelfeed/I_28  ( .A(\pixelfeed/N225 ), .Z(\pixelfeed/N226 ) );
  GTECH_AND2 \pixelfeed/C701  ( .A(\pixelfeed/N212 ), .B(\pixelfeed/N224 ), 
        .Z(\pixelfeed/N225 ) );
  GTECH_AND2 \pixelfeed/C700  ( .A(fml_stb), .B(\pixelfeed/N151 ), .Z(
        \pixelfeed/N224 ) );
  GTECH_NOT \pixelfeed/I_27  ( .A(\pixelfeed/N222 ), .Z(\pixelfeed/N223 ) );
  GTECH_OR2 \pixelfeed/C698  ( .A(\pixelfeed/N203 ), .B(\pixelfeed/N221 ), .Z(
        \pixelfeed/N222 ) );
  GTECH_OR2 \pixelfeed/C697  ( .A(\pixelfeed/N199 ), .B(\pixelfeed/N220 ), .Z(
        \pixelfeed/N221 ) );
  GTECH_OR2 \pixelfeed/C696  ( .A(\pixelfeed/N195 ), .B(\pixelfeed/N219 ), .Z(
        \pixelfeed/N220 ) );
  GTECH_OR2 \pixelfeed/C695  ( .A(fml_stb), .B(\pixelfeed/N218 ), .Z(
        \pixelfeed/N219 ) );
  GTECH_OR2 \pixelfeed/C694  ( .A(\pixelfeed/N187 ), .B(\pixelfeed/N217 ), .Z(
        \pixelfeed/N218 ) );
  GTECH_OR2 \pixelfeed/C693  ( .A(\pixelfeed/N183 ), .B(\pixelfeed/N216 ), .Z(
        \pixelfeed/N217 ) );
  GTECH_OR2 \pixelfeed/C692  ( .A(\pixelfeed/N179 ), .B(\pixelfeed/N215 ), .Z(
        \pixelfeed/N216 ) );
  GTECH_OR2 \pixelfeed/C691  ( .A(\pixelfeed/N175 ), .B(\pixelfeed/N214 ), .Z(
        \pixelfeed/N215 ) );
  GTECH_OR2 \pixelfeed/C690  ( .A(\pixelfeed/N171 ), .B(\pixelfeed/N167 ), .Z(
        \pixelfeed/N214 ) );
  GTECH_NOT \pixelfeed/I_26  ( .A(fml_ack), .Z(\pixelfeed/N212 ) );
  GTECH_NOT \pixelfeed/I_25  ( .A(dcb_hit), .Z(\pixelfeed/N210 ) );
  GTECH_NOT \pixelfeed/I_24  ( .A(\pixelfeed/N204 ), .Z(\pixelfeed/N205 ) );
  GTECH_NOT \pixelfeed/I_23  ( .A(vga_rst), .Z(\pixelfeed/N266 ) );
  GTECH_NOT \pixelfeed/I_22  ( .A(pixel_valid), .Z(\pixelfeed/N265 ) );
  GTECH_AND2 \pixelfeed/C678  ( .A(\pixelfeed/N265 ), .B(\pixelfeed/N266 ), 
        .Z(\pixelfeed/N204 ) );
  GTECH_BUF \pixelfeed/B_40  ( .A(\pixelfeed/N191 ), .Z(fml_stb) );
  GTECH_NOT \pixelfeed/I_21  ( .A(\pixelfeed/N202 ), .Z(\pixelfeed/N203 ) );
  GTECH_NOT \pixelfeed/I_20  ( .A(\pixelfeed/N198 ), .Z(\pixelfeed/N199 ) );
  GTECH_NOT \pixelfeed/I_19  ( .A(\pixelfeed/N194 ), .Z(\pixelfeed/N195 ) );
  GTECH_NOT \pixelfeed/I_18  ( .A(\pixelfeed/N190 ), .Z(\pixelfeed/N191 ) );
  GTECH_NOT \pixelfeed/I_17  ( .A(\pixelfeed/N186 ), .Z(\pixelfeed/N187 ) );
  GTECH_NOT \pixelfeed/I_16  ( .A(\pixelfeed/N182 ), .Z(\pixelfeed/N183 ) );
  GTECH_NOT \pixelfeed/I_15  ( .A(\pixelfeed/N178 ), .Z(\pixelfeed/N179 ) );
  GTECH_NOT \pixelfeed/I_14  ( .A(\pixelfeed/N174 ), .Z(\pixelfeed/N175 ) );
  GTECH_NOT \pixelfeed/I_13  ( .A(\pixelfeed/N170 ), .Z(\pixelfeed/N171 ) );
  GTECH_NOT \pixelfeed/I_12  ( .A(\pixelfeed/state[0] ), .Z(\pixelfeed/N164 )
         );
  GTECH_NOT \pixelfeed/I_11  ( .A(\pixelfeed/state[1] ), .Z(\pixelfeed/N163 )
         );
  GTECH_NOT \pixelfeed/I_10  ( .A(\pixelfeed/state[2] ), .Z(\pixelfeed/N162 )
         );
  GTECH_NOT \pixelfeed/I_9  ( .A(\pixelfeed/state[3] ), .Z(\pixelfeed/N161 )
         );
  GTECH_NOT \pixelfeed/I_8  ( .A(\pixelfeed/ignore ), .Z(\pixelfeed/N160 ) );
  GTECH_AND2 \pixelfeed/C638  ( .A(\pixelfeed/ignore_clear ), .B(
        \pixelfeed/N158 ), .Z(\pixelfeed/N159 ) );
  GTECH_NOT \pixelfeed/I_7  ( .A(\pixelfeed/N157 ), .Z(\pixelfeed/N158 ) );
  GTECH_BUF \pixelfeed/B_39  ( .A(vga_rst), .Z(\pixelfeed/N157 ) );
  GTECH_NOT \pixelfeed/I_6  ( .A(sys_rst), .Z(\pixelfeed/N151 ) );
  GTECH_BUF \pixelfeed/B_38  ( .A(dcb_stb), .Z() );
  GTECH_NOT \pixelfeed/I_5  ( .A(dcb_stb), .Z(\pixelfeed/N146 ) );
  GTECH_AND2 \pixelfeed/C627  ( .A(\pixelfeed/ignore_clear ), .B(
        \pixelfeed/N144 ), .Z(\pixelfeed/N145 ) );
  GTECH_NOT \pixelfeed/I_4  ( .A(sys_rst), .Z(\pixelfeed/N144 ) );
  GTECH_AND2 \pixelfeed/C625  ( .A(\pixelfeed/N63 ), .B(\pixelfeed/N64 ), .Z()
         );
  GTECH_NOT \pixelfeed/I_3  ( .A(\pixelfeed/sof ), .Z(\pixelfeed/N64 ) );
  GTECH_BUF \pixelfeed/B_37  ( .A(\pixelfeed/N145 ), .Z(\pixelfeed/N63 ) );
  GTECH_AND2 \pixelfeed/C619  ( .A(\pixelfeed/sof ), .B(
        \pixelfeed/ignore_clear ), .Z(baseaddress_ack) );
  GTECH_AND2 \pixelfeed/C618  ( .A(\pixelfeed/N37 ), .B(\pixelfeed/N61 ), .Z()
         );
  GTECH_AND2 \pixelfeed/C617  ( .A(\pixelfeed/ignore_clear ), .B(
        \pixelfeed/N61 ), .Z(\pixelfeed/N62 ) );
  GTECH_NOT \pixelfeed/I_2  ( .A(\pixelfeed/N36 ), .Z(\pixelfeed/N61 ) );
  GTECH_AND2 \pixelfeed/C615  ( .A(\pixelfeed/N37 ), .B(\pixelfeed/N39 ), .Z(
        \pixelfeed/N40 ) );
  GTECH_NOT \pixelfeed/I_1  ( .A(\pixelfeed/N38 ), .Z(\pixelfeed/N39 ) );
  GTECH_BUF \pixelfeed/B_36  ( .A(\pixelfeed/N62 ), .Z(\pixelfeed/N37 ) );
  GTECH_BUF \pixelfeed/B_35  ( .A(vga_rst), .Z(\pixelfeed/N36 ) );
  GTECH_NOT \pixelfeed/I_0  ( .A(\pixelfeed/fifo_source_cache ), .Z(
        \pixelfeed/N35 ) );
  MULT_UNS_OP \pixelfeed/mult_add_84_aco  ( .A({\pixelfeed/bcounter[17] , 
        \pixelfeed/bcounter[16] , \pixelfeed/bcounter[15] , 
        \pixelfeed/bcounter[14] , \pixelfeed/bcounter[13] , 
        \pixelfeed/bcounter[12] , \pixelfeed/bcounter[11] , 
        \pixelfeed/bcounter[10] , \pixelfeed/bcounter[9] , 
        \pixelfeed/bcounter[8] , \pixelfeed/bcounter[7] , 
        \pixelfeed/bcounter[6] , \pixelfeed/bcounter[5] , 
        \pixelfeed/bcounter[4] , \pixelfeed/bcounter[3] , 
        \pixelfeed/bcounter[2] , \pixelfeed/bcounter[1] , 
        \pixelfeed/bcounter[0] }), .B(\pixelfeed/N246 ), .Z({\pixelfeed/N264 , 
        \pixelfeed/N263 , \pixelfeed/N262 , \pixelfeed/N261 , \pixelfeed/N260 , 
        \pixelfeed/N259 , \pixelfeed/N258 , \pixelfeed/N257 , \pixelfeed/N256 , 
        \pixelfeed/N255 , \pixelfeed/N254 , \pixelfeed/N253 , \pixelfeed/N252 , 
        \pixelfeed/N251 , \pixelfeed/N250 , \pixelfeed/N249 , \pixelfeed/N248 , 
        \pixelfeed/N247 }) );
  GTECH_BUF \pixelfeed/B_34  ( .A(\pixelfeed/N203 ), .Z(\pixelfeed/N34 ) );
  GTECH_BUF \pixelfeed/B_33  ( .A(\pixelfeed/N199 ), .Z(\pixelfeed/N33 ) );
  GTECH_BUF \pixelfeed/B_32  ( .A(\pixelfeed/N195 ), .Z(\pixelfeed/N32 ) );
  GTECH_BUF \pixelfeed/B_31  ( .A(fml_stb), .Z(\pixelfeed/N31 ) );
  GTECH_BUF \pixelfeed/B_30  ( .A(\pixelfeed/N187 ), .Z(\pixelfeed/N30 ) );
  GTECH_BUF \pixelfeed/B_29  ( .A(\pixelfeed/N183 ), .Z(\pixelfeed/N29 ) );
  GTECH_BUF \pixelfeed/B_28  ( .A(\pixelfeed/N179 ), .Z(\pixelfeed/N28 ) );
  GTECH_BUF \pixelfeed/B_27  ( .A(\pixelfeed/N244 ), .Z(\pixelfeed/N27 ) );
  SELECT_OP \pixelfeed/C600  ( .DATA1(1'b0), .DATA2(\pixelfeed/N211 ), .DATA3(
        \pixelfeed/N160 ), .DATA4(\pixelfeed/N160 ), .DATA5(\pixelfeed/N160 ), 
        .DATA6(\pixelfeed/N213 ), .DATA7(\pixelfeed/N160 ), .DATA8(
        \pixelfeed/N160 ), .DATA9(\pixelfeed/N160 ), .CONTROL1(\pixelfeed/N27 ), .CONTROL2(\pixelfeed/N16 ), .CONTROL3(\pixelfeed/N28 ), .CONTROL4(
        \pixelfeed/N29 ), .CONTROL5(\pixelfeed/N30 ), .CONTROL6(
        \pixelfeed/N31 ), .CONTROL7(\pixelfeed/N32 ), .CONTROL8(
        \pixelfeed/N33 ), .CONTROL9(\pixelfeed/N34 ), .Z(\pixelfeed/fifo_stb )
         );
  GTECH_BUF \pixelfeed/B_26  ( .A(\pixelfeed/N243 ), .Z(\pixelfeed/N26 ) );
  GTECH_BUF \pixelfeed/B_25  ( .A(\pixelfeed/N242 ), .Z(\pixelfeed/N25 ) );
  SELECT_OP \pixelfeed/C599  ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(dcb_hit), 
        .CONTROL1(\pixelfeed/N25 ), .CONTROL2(\pixelfeed/N26 ), .CONTROL3(
        \pixelfeed/N16 ), .Z(dcb_stb) );
  GTECH_BUF \pixelfeed/B_24  ( .A(\pixelfeed/N239 ), .Z(\pixelfeed/N24 ) );
  SELECT_OP \pixelfeed/C598  ( .DATA1(\pixelfeed/N204 ), .DATA2(1'b0), 
        .CONTROL1(\pixelfeed/N14 ), .CONTROL2(\pixelfeed/N24 ), .Z(
        \pixelfeed/ignore_clear ) );
  GTECH_BUF \pixelfeed/B_23  ( .A(\pixelfeed/N237 ), .Z(\pixelfeed/N23 ) );
  GTECH_BUF \pixelfeed/B_22  ( .A(\pixelfeed/N236 ), .Z(\pixelfeed/N22 ) );
  SELECT_OP \pixelfeed/C597  ( .DATA1(\pixelfeed/N209 ), .DATA2(1'b0), .DATA3(
        1'b1), .DATA4(\pixelfeed/state[3] ), .CONTROL1(\pixelfeed/N14 ), 
        .CONTROL2(\pixelfeed/N22 ), .CONTROL3(\pixelfeed/N23 ), .CONTROL4(
        \pixelfeed/N223 ), .Z(\pixelfeed/next_state [3]) );
  GTECH_BUF \pixelfeed/B_21  ( .A(\pixelfeed/N233 ), .Z(\pixelfeed/N21 ) );
  GTECH_BUF \pixelfeed/B_20  ( .A(\pixelfeed/N232 ), .Z(\pixelfeed/N20 ) );
  SELECT_OP \pixelfeed/C596  ( .DATA1(\pixelfeed/N208 ), .DATA2(1'b0), .DATA3(
        \pixelfeed/N210 ), .DATA4(1'b1), .DATA5(\pixelfeed/state[2] ), 
        .CONTROL1(\pixelfeed/N14 ), .CONTROL2(\pixelfeed/N20 ), .CONTROL3(
        \pixelfeed/N16 ), .CONTROL4(\pixelfeed/N21 ), .CONTROL5(
        \pixelfeed/N223 ), .Z(\pixelfeed/next_state [2]) );
  GTECH_BUF \pixelfeed/B_19  ( .A(\pixelfeed/N231 ), .Z(\pixelfeed/N19 ) );
  GTECH_BUF \pixelfeed/B_18  ( .A(\pixelfeed/N229 ), .Z(\pixelfeed/N18 ) );
  SELECT_OP \pixelfeed/C595  ( .DATA1(\pixelfeed/N207 ), .DATA2(1'b1), .DATA3(
        1'b0), .DATA4(\pixelfeed/state[1] ), .CONTROL1(\pixelfeed/N14 ), 
        .CONTROL2(\pixelfeed/N18 ), .CONTROL3(\pixelfeed/N19 ), .CONTROL4(
        \pixelfeed/N223 ), .Z(\pixelfeed/next_state [1]) );
  GTECH_BUF \pixelfeed/B_17  ( .A(\pixelfeed/N228 ), .Z(\pixelfeed/N17 ) );
  GTECH_BUF \pixelfeed/B_16  ( .A(\pixelfeed/N175 ), .Z(\pixelfeed/N16 ) );
  GTECH_BUF \pixelfeed/B_15  ( .A(\pixelfeed/N227 ), .Z(\pixelfeed/N15 ) );
  GTECH_BUF \pixelfeed/B_14  ( .A(\pixelfeed/N167 ), .Z(\pixelfeed/N14 ) );
  SELECT_OP \pixelfeed/C594  ( .DATA1(\pixelfeed/N206 ), .DATA2(1'b0), .DATA3(
        dcb_hit), .DATA4(1'b1), .DATA5(\pixelfeed/state[0] ), .CONTROL1(
        \pixelfeed/N14 ), .CONTROL2(\pixelfeed/N15 ), .CONTROL3(
        \pixelfeed/N16 ), .CONTROL4(\pixelfeed/N17 ), .CONTROL5(
        \pixelfeed/N223 ), .Z(\pixelfeed/next_state [0]) );
  GTECH_BUF \pixelfeed/B_13  ( .A(\pixelfeed/N212 ), .Z(\pixelfeed/N13 ) );
  GTECH_BUF \pixelfeed/B_12  ( .A(fml_ack), .Z(\pixelfeed/N12 ) );
  SELECT_OP \pixelfeed/C593  ( .DATA1(\pixelfeed/N160 ), .DATA2(1'b0), 
        .CONTROL1(\pixelfeed/N12 ), .CONTROL2(\pixelfeed/N13 ), .Z(
        \pixelfeed/N213 ) );
  GTECH_BUF \pixelfeed/B_11  ( .A(\pixelfeed/N210 ), .Z(\pixelfeed/N11 ) );
  GTECH_BUF \pixelfeed/B_10  ( .A(dcb_hit), .Z(\pixelfeed/N10 ) );
  SELECT_OP \pixelfeed/C592  ( .DATA1(\pixelfeed/N160 ), .DATA2(1'b0), 
        .CONTROL1(\pixelfeed/N10 ), .CONTROL2(\pixelfeed/N11 ), .Z(
        \pixelfeed/N211 ) );
  GTECH_BUF \pixelfeed/B_9  ( .A(\pixelfeed/N204 ), .Z(\pixelfeed/N9 ) );
  SELECT_OP \pixelfeed/C591  ( .DATA1({1'b0, 1'b0, 1'b0, 1'b1}), .DATA2({
        \pixelfeed/state[3] , \pixelfeed/state[2] , \pixelfeed/state[1] , 
        \pixelfeed/state[0] }), .CONTROL1(\pixelfeed/N9 ), .CONTROL2(
        \pixelfeed/N205 ), .Z({\pixelfeed/N209 , \pixelfeed/N208 , 
        \pixelfeed/N207 , \pixelfeed/N206 }) );
  GTECH_BUF \pixelfeed/B_8  ( .A(\pixelfeed/N151 ), .Z(\pixelfeed/N8 ) );
  SELECT_OP \pixelfeed/C590  ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0}), .DATA2(
        \pixelfeed/next_state ), .CONTROL1(\pixelfeed/N5 ), .CONTROL2(
        \pixelfeed/N8 ), .Z({\pixelfeed/N155 , \pixelfeed/N154 , 
        \pixelfeed/N153 , \pixelfeed/N152 }) );
  GTECH_BUF \pixelfeed/B_7  ( .A(\pixelfeed/N146 ), .Z(\pixelfeed/N7 ) );
  GTECH_BUF \pixelfeed/B_6  ( .A(dcb_stb), .Z(\pixelfeed/N6 ) );
  SELECT_OP \pixelfeed/C589  ( .DATA1({\pixelfeed/N148 , \pixelfeed/N147 }), 
        .DATA2({1'b0, 1'b0}), .CONTROL1(\pixelfeed/N6 ), .CONTROL2(
        \pixelfeed/N7 ), .Z({\pixelfeed/N150 , \pixelfeed/N149 }) );
  GTECH_BUF \pixelfeed/B_5  ( .A(sys_rst), .Z(\pixelfeed/N5 ) );
  SELECT_OP \pixelfeed/C588  ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .DATA2({
        \pixelfeed/N116 , \pixelfeed/N115 , \pixelfeed/N114 , \pixelfeed/N113 , 
        \pixelfeed/N112 , \pixelfeed/N111 , \pixelfeed/N110 , \pixelfeed/N109 , 
        \pixelfeed/N108 , \pixelfeed/N107 , \pixelfeed/N106 , \pixelfeed/N105 , 
        \pixelfeed/N104 , \pixelfeed/N103 , \pixelfeed/N102 , \pixelfeed/N101 , 
        \pixelfeed/N100 , \pixelfeed/N99 , \pixelfeed/N98 , \pixelfeed/N97 , 
        \pixelfeed/N96 , \pixelfeed/N95 , \pixelfeed/N94 , \pixelfeed/N93 , 
        \pixelfeed/N92 , \pixelfeed/N91 }), .CONTROL1(\pixelfeed/N5 ), 
        .CONTROL2(\pixelfeed/N145 ), .Z({\pixelfeed/N143 , \pixelfeed/N142 , 
        \pixelfeed/N141 , \pixelfeed/N140 , \pixelfeed/N139 , \pixelfeed/N138 , 
        \pixelfeed/N137 , \pixelfeed/N136 , \pixelfeed/N135 , \pixelfeed/N134 , 
        \pixelfeed/N133 , \pixelfeed/N132 , \pixelfeed/N131 , \pixelfeed/N130 , 
        \pixelfeed/N129 , \pixelfeed/N128 , \pixelfeed/N127 , \pixelfeed/N126 , 
        \pixelfeed/N125 , \pixelfeed/N124 , \pixelfeed/N123 , \pixelfeed/N122 , 
        \pixelfeed/N121 , \pixelfeed/N120 , \pixelfeed/N119 , \pixelfeed/N118 }) );
  GTECH_BUF \pixelfeed/B_4  ( .A(\pixelfeed/N64 ), .Z(\pixelfeed/N4 ) );
  GTECH_BUF \pixelfeed/B_3  ( .A(\pixelfeed/sof ), .Z(\pixelfeed/N3 ) );
  SELECT_OP \pixelfeed/C587  ( .DATA1(baseaddress), .DATA2({\pixelfeed/N90 , 
        \pixelfeed/N89 , \pixelfeed/N88 , \pixelfeed/N87 , \pixelfeed/N86 , 
        \pixelfeed/N85 , \pixelfeed/N84 , \pixelfeed/N83 , \pixelfeed/N82 , 
        \pixelfeed/N81 , \pixelfeed/N80 , \pixelfeed/N79 , \pixelfeed/N78 , 
        \pixelfeed/N77 , \pixelfeed/N76 , \pixelfeed/N75 , \pixelfeed/N74 , 
        \pixelfeed/N73 , \pixelfeed/N72 , \pixelfeed/N71 , \pixelfeed/N70 , 
        \pixelfeed/N69 , \pixelfeed/N68 , \pixelfeed/N67 , \pixelfeed/N66 , 
        \pixelfeed/N65 }), .CONTROL1(\pixelfeed/N3 ), .CONTROL2(\pixelfeed/N4 ), .Z({\pixelfeed/N116 , \pixelfeed/N115 , \pixelfeed/N114 , \pixelfeed/N113 , 
        \pixelfeed/N112 , \pixelfeed/N111 , \pixelfeed/N110 , \pixelfeed/N109 , 
        \pixelfeed/N108 , \pixelfeed/N107 , \pixelfeed/N106 , \pixelfeed/N105 , 
        \pixelfeed/N104 , \pixelfeed/N103 , \pixelfeed/N102 , \pixelfeed/N101 , 
        \pixelfeed/N100 , \pixelfeed/N99 , \pixelfeed/N98 , \pixelfeed/N97 , 
        \pixelfeed/N96 , \pixelfeed/N95 , \pixelfeed/N94 , \pixelfeed/N93 , 
        \pixelfeed/N92 , \pixelfeed/N91 }) );
  GTECH_BUF \pixelfeed/B_2  ( .A(\pixelfeed/N36 ), .Z(\pixelfeed/N2 ) );
  SELECT_OP \pixelfeed/C586  ( .DATA1(1'b1), .DATA2(\pixelfeed/N38 ), 
        .CONTROL1(\pixelfeed/N2 ), .CONTROL2(\pixelfeed/N62 ), .Z(
        \pixelfeed/N60 ) );
  GTECH_BUF \pixelfeed/B_1  ( .A(\pixelfeed/N35 ), .Z(\pixelfeed/N1 ) );
  GTECH_BUF \pixelfeed/B_0  ( .A(\pixelfeed/fifo_source_cache ), .Z(
        \pixelfeed/N0 ) );
  SELECT_OP \pixelfeed/C583  ( .DATA1(dcb_dat), .DATA2(fml_di), .CONTROL1(
        \pixelfeed/N0 ), .CONTROL2(\pixelfeed/N1 ), .Z({
        \pixelfeed/n_0_net__63_ , \pixelfeed/n_0_net__62_ , 
        \pixelfeed/n_0_net__61_ , \pixelfeed/n_0_net__60_ , 
        \pixelfeed/n_0_net__59_ , \pixelfeed/n_0_net__58_ , 
        \pixelfeed/n_0_net__57_ , \pixelfeed/n_0_net__56_ , 
        \pixelfeed/n_0_net__55_ , \pixelfeed/n_0_net__54_ , 
        \pixelfeed/n_0_net__53_ , \pixelfeed/n_0_net__52_ , 
        \pixelfeed/n_0_net__51_ , \pixelfeed/n_0_net__50_ , 
        \pixelfeed/n_0_net__49_ , \pixelfeed/n_0_net__48_ , 
        \pixelfeed/n_0_net__47_ , \pixelfeed/n_0_net__46_ , 
        \pixelfeed/n_0_net__45_ , \pixelfeed/n_0_net__44_ , 
        \pixelfeed/n_0_net__43_ , \pixelfeed/n_0_net__42_ , 
        \pixelfeed/n_0_net__41_ , \pixelfeed/n_0_net__40_ , 
        \pixelfeed/n_0_net__39_ , \pixelfeed/n_0_net__38_ , 
        \pixelfeed/n_0_net__37_ , \pixelfeed/n_0_net__36_ , 
        \pixelfeed/n_0_net__35_ , \pixelfeed/n_0_net__34_ , 
        \pixelfeed/n_0_net__33_ , \pixelfeed/n_0_net__32_ , 
        \pixelfeed/n_0_net__31_ , \pixelfeed/n_0_net__30_ , 
        \pixelfeed/n_0_net__29_ , \pixelfeed/n_0_net__28_ , 
        \pixelfeed/n_0_net__27_ , \pixelfeed/n_0_net__26_ , 
        \pixelfeed/n_0_net__25_ , \pixelfeed/n_0_net__24_ , 
        \pixelfeed/n_0_net__23_ , \pixelfeed/n_0_net__22_ , 
        \pixelfeed/n_0_net__21_ , \pixelfeed/n_0_net__20_ , 
        \pixelfeed/n_0_net__19_ , \pixelfeed/n_0_net__18_ , 
        \pixelfeed/n_0_net__17_ , \pixelfeed/n_0_net__16_ , 
        \pixelfeed/n_0_net__15_ , \pixelfeed/n_0_net__14_ , 
        \pixelfeed/n_0_net__13_ , \pixelfeed/n_0_net__12_ , 
        \pixelfeed/n_0_net__11_ , \pixelfeed/n_0_net__10_ , 
        \pixelfeed/n_0_net__9_ , \pixelfeed/n_0_net__8_ , 
        \pixelfeed/n_0_net__7_ , \pixelfeed/n_0_net__6_ , 
        \pixelfeed/n_0_net__5_ , \pixelfeed/n_0_net__4_ , 
        \pixelfeed/n_0_net__3_ , \pixelfeed/n_0_net__2_ , 
        \pixelfeed/n_0_net__1_ , \pixelfeed/n_0_net__0_ }) );
  ADD_UNS_OP \pixelfeed/add_84_aco  ( .A({\pixelfeed/N264 , \pixelfeed/N263 , 
        \pixelfeed/N262 , \pixelfeed/N261 , \pixelfeed/N260 , \pixelfeed/N259 , 
        \pixelfeed/N258 , \pixelfeed/N257 , \pixelfeed/N256 , \pixelfeed/N255 , 
        \pixelfeed/N254 , \pixelfeed/N253 , \pixelfeed/N252 , \pixelfeed/N251 , 
        \pixelfeed/N250 , \pixelfeed/N249 , \pixelfeed/N248 , \pixelfeed/N247 }), .B(1'b1), .Z({\pixelfeed/N59 , \pixelfeed/N58 , \pixelfeed/N57 , 
        \pixelfeed/N56 , \pixelfeed/N55 , \pixelfeed/N54 , \pixelfeed/N53 , 
        \pixelfeed/N52 , \pixelfeed/N51 , \pixelfeed/N50 , \pixelfeed/N49 , 
        \pixelfeed/N48 , \pixelfeed/N47 , \pixelfeed/N46 , \pixelfeed/N45 , 
        \pixelfeed/N44 , \pixelfeed/N43 , \pixelfeed/N42 }) );
  ADD_UNS_OP \pixelfeed/add_104  ( .A(fml_adr), .B({1'b1, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .Z({\pixelfeed/N90 , \pixelfeed/N89 , \pixelfeed/N88 , 
        \pixelfeed/N87 , \pixelfeed/N86 , \pixelfeed/N85 , \pixelfeed/N84 , 
        \pixelfeed/N83 , \pixelfeed/N82 , \pixelfeed/N81 , \pixelfeed/N80 , 
        \pixelfeed/N79 , \pixelfeed/N78 , \pixelfeed/N77 , \pixelfeed/N76 , 
        \pixelfeed/N75 , \pixelfeed/N74 , \pixelfeed/N73 , \pixelfeed/N72 , 
        \pixelfeed/N71 , \pixelfeed/N70 , \pixelfeed/N69 , \pixelfeed/N68 , 
        \pixelfeed/N67 , \pixelfeed/N66 , \pixelfeed/N65 }) );
  GTECH_OR2 \pixelfeed/C531  ( .A(sys_rst), .B(\pixelfeed/N145 ), .Z(
        \pixelfeed/N117 ) );
  GTECH_OR2 \pixelfeed/C493  ( .A(\pixelfeed/N36 ), .B(\pixelfeed/N62 ), .Z(
        \pixelfeed/N41 ) );
  GTECH_OR2 \pixelfeed/C491  ( .A(\pixelfeed/N157 ), .B(\pixelfeed/N159 ), .Z(
        \pixelfeed/N156 ) );
  ADD_UNS_OP \pixelfeed/add_114  ( .A(dcb_adr[4:3]), .B(1'b1), .Z({
        \pixelfeed/N148 , \pixelfeed/N147 }) );
  GTECH_OR3 \pixelfeed/C485  ( .A(\pixelfeed/N167 ), .B(\pixelfeed/N171 ), .C(
        \pixelfeed/N223 ), .Z(\pixelfeed/N244 ) );
  GTECH_OR4 \pixelfeed/C483  ( .A(\pixelfeed/N175 ), .B(\pixelfeed/N179 ), .C(
        \pixelfeed/N183 ), .D(\pixelfeed/N187 ), .Z(
        \pixelfeed/fifo_source_cache ) );
  GTECH_OR3 \pixelfeed/C478  ( .A(\pixelfeed/N171 ), .B(\pixelfeed/N179 ), .C(
        \pixelfeed/N183 ), .Z(\pixelfeed/N243 ) );
  GTECH_OR2 \pixelfeed/C477  ( .A(\pixelfeed/N240 ), .B(\pixelfeed/N241 ), .Z(
        \pixelfeed/N242 ) );
  GTECH_OR2 \pixelfeed/C476  ( .A(\pixelfeed/N203 ), .B(\pixelfeed/N223 ), .Z(
        \pixelfeed/N241 ) );
  GTECH_OR5 \pixelfeed/C475  ( .A(\pixelfeed/N167 ), .B(\pixelfeed/N187 ), .C(
        fml_stb), .D(\pixelfeed/N195 ), .E(\pixelfeed/N199 ), .Z(
        \pixelfeed/N240 ) );
  GTECH_OR2 \pixelfeed/C473  ( .A(\pixelfeed/N234 ), .B(\pixelfeed/N238 ), .Z(
        \pixelfeed/N239 ) );
  GTECH_OR5 \pixelfeed/C472  ( .A(fml_stb), .B(\pixelfeed/N195 ), .C(
        \pixelfeed/N199 ), .D(\pixelfeed/N203 ), .E(\pixelfeed/N223 ), .Z(
        \pixelfeed/N238 ) );
  GTECH_OR2 \pixelfeed/C469  ( .A(\pixelfeed/N195 ), .B(\pixelfeed/N199 ), .Z(
        \pixelfeed/N237 ) );
  GTECH_OR2 \pixelfeed/C468  ( .A(\pixelfeed/N234 ), .B(\pixelfeed/N235 ), .Z(
        \pixelfeed/N236 ) );
  GTECH_OR2 \pixelfeed/C467  ( .A(fml_stb), .B(\pixelfeed/N203 ), .Z(
        \pixelfeed/N235 ) );
  GTECH_OR5 \pixelfeed/C466  ( .A(\pixelfeed/N171 ), .B(\pixelfeed/N175 ), .C(
        \pixelfeed/N179 ), .D(\pixelfeed/N183 ), .E(\pixelfeed/N187 ), .Z(
        \pixelfeed/N234 ) );
  GTECH_OR3 \pixelfeed/C464  ( .A(\pixelfeed/N179 ), .B(\pixelfeed/N183 ), .C(
        fml_stb), .Z(\pixelfeed/N233 ) );
  GTECH_OR5 \pixelfeed/C463  ( .A(\pixelfeed/N171 ), .B(\pixelfeed/N187 ), .C(
        \pixelfeed/N195 ), .D(\pixelfeed/N199 ), .E(\pixelfeed/N203 ), .Z(
        \pixelfeed/N232 ) );
  GTECH_OR2 \pixelfeed/C461  ( .A(\pixelfeed/N230 ), .B(\pixelfeed/N203 ), .Z(
        \pixelfeed/N231 ) );
  GTECH_OR5 \pixelfeed/C460  ( .A(\pixelfeed/N179 ), .B(\pixelfeed/N183 ), .C(
        \pixelfeed/N187 ), .D(\pixelfeed/N195 ), .E(\pixelfeed/N199 ), .Z(
        \pixelfeed/N230 ) );
  GTECH_OR3 \pixelfeed/C459  ( .A(\pixelfeed/N171 ), .B(\pixelfeed/N175 ), .C(
        fml_stb), .Z(\pixelfeed/N229 ) );
  GTECH_OR3 \pixelfeed/C457  ( .A(\pixelfeed/N183 ), .B(fml_stb), .C(
        \pixelfeed/N199 ), .Z(\pixelfeed/N228 ) );
  GTECH_OR5 \pixelfeed/C456  ( .A(\pixelfeed/N171 ), .B(\pixelfeed/N179 ), .C(
        \pixelfeed/N187 ), .D(\pixelfeed/N195 ), .E(\pixelfeed/N203 ), .Z(
        \pixelfeed/N227 ) );
  GTECH_OR2 \pixelfeed/C332  ( .A(\pixelfeed/N200 ), .B(\pixelfeed/N201 ), .Z(
        \pixelfeed/N202 ) );
  GTECH_OR2 \pixelfeed/C331  ( .A(\pixelfeed/state[1] ), .B(\pixelfeed/N164 ), 
        .Z(\pixelfeed/N201 ) );
  GTECH_OR2 \pixelfeed/C330  ( .A(\pixelfeed/N161 ), .B(\pixelfeed/state[2] ), 
        .Z(\pixelfeed/N200 ) );
  GTECH_OR2 \pixelfeed/C326  ( .A(\pixelfeed/N196 ), .B(\pixelfeed/N197 ), .Z(
        \pixelfeed/N198 ) );
  GTECH_OR2 \pixelfeed/C325  ( .A(\pixelfeed/state[1] ), .B(
        \pixelfeed/state[0] ), .Z(\pixelfeed/N197 ) );
  GTECH_OR2 \pixelfeed/C324  ( .A(\pixelfeed/N161 ), .B(\pixelfeed/state[2] ), 
        .Z(\pixelfeed/N196 ) );
  GTECH_OR2 \pixelfeed/C321  ( .A(\pixelfeed/N192 ), .B(\pixelfeed/N193 ), .Z(
        \pixelfeed/N194 ) );
  GTECH_OR2 \pixelfeed/C320  ( .A(\pixelfeed/N163 ), .B(\pixelfeed/N164 ), .Z(
        \pixelfeed/N193 ) );
  GTECH_OR2 \pixelfeed/C319  ( .A(\pixelfeed/state[3] ), .B(\pixelfeed/N162 ), 
        .Z(\pixelfeed/N192 ) );
  GTECH_OR2 \pixelfeed/C314  ( .A(\pixelfeed/N188 ), .B(\pixelfeed/N189 ), .Z(
        \pixelfeed/N190 ) );
  GTECH_OR2 \pixelfeed/C313  ( .A(\pixelfeed/N163 ), .B(\pixelfeed/state[0] ), 
        .Z(\pixelfeed/N189 ) );
  GTECH_OR2 \pixelfeed/C312  ( .A(\pixelfeed/state[3] ), .B(\pixelfeed/N162 ), 
        .Z(\pixelfeed/N188 ) );
  GTECH_OR2 \pixelfeed/C308  ( .A(\pixelfeed/N184 ), .B(\pixelfeed/N185 ), .Z(
        \pixelfeed/N186 ) );
  GTECH_OR2 \pixelfeed/C307  ( .A(\pixelfeed/state[1] ), .B(\pixelfeed/N164 ), 
        .Z(\pixelfeed/N185 ) );
  GTECH_OR2 \pixelfeed/C306  ( .A(\pixelfeed/state[3] ), .B(\pixelfeed/N162 ), 
        .Z(\pixelfeed/N184 ) );
  GTECH_OR2 \pixelfeed/C302  ( .A(\pixelfeed/N180 ), .B(\pixelfeed/N181 ), .Z(
        \pixelfeed/N182 ) );
  GTECH_OR2 \pixelfeed/C301  ( .A(\pixelfeed/state[1] ), .B(
        \pixelfeed/state[0] ), .Z(\pixelfeed/N181 ) );
  GTECH_OR2 \pixelfeed/C300  ( .A(\pixelfeed/state[3] ), .B(\pixelfeed/N162 ), 
        .Z(\pixelfeed/N180 ) );
  GTECH_OR2 \pixelfeed/C297  ( .A(\pixelfeed/N176 ), .B(\pixelfeed/N177 ), .Z(
        \pixelfeed/N178 ) );
  GTECH_OR2 \pixelfeed/C296  ( .A(\pixelfeed/N163 ), .B(\pixelfeed/N164 ), .Z(
        \pixelfeed/N177 ) );
  GTECH_OR2 \pixelfeed/C295  ( .A(\pixelfeed/state[3] ), .B(
        \pixelfeed/state[2] ), .Z(\pixelfeed/N176 ) );
  GTECH_OR2 \pixelfeed/C291  ( .A(\pixelfeed/N172 ), .B(\pixelfeed/N173 ), .Z(
        \pixelfeed/N174 ) );
  GTECH_OR2 \pixelfeed/C290  ( .A(\pixelfeed/N163 ), .B(\pixelfeed/state[0] ), 
        .Z(\pixelfeed/N173 ) );
  GTECH_OR2 \pixelfeed/C289  ( .A(\pixelfeed/state[3] ), .B(
        \pixelfeed/state[2] ), .Z(\pixelfeed/N172 ) );
  GTECH_OR2 \pixelfeed/C286  ( .A(\pixelfeed/N168 ), .B(\pixelfeed/N169 ), .Z(
        \pixelfeed/N170 ) );
  GTECH_OR2 \pixelfeed/C285  ( .A(\pixelfeed/state[1] ), .B(\pixelfeed/N164 ), 
        .Z(\pixelfeed/N169 ) );
  GTECH_OR2 \pixelfeed/C284  ( .A(\pixelfeed/state[3] ), .B(
        \pixelfeed/state[2] ), .Z(\pixelfeed/N168 ) );
  GTECH_AND2 \pixelfeed/C282  ( .A(\pixelfeed/N165 ), .B(\pixelfeed/N166 ), 
        .Z(\pixelfeed/N167 ) );
  GTECH_AND2 \pixelfeed/C281  ( .A(\pixelfeed/N163 ), .B(\pixelfeed/N164 ), 
        .Z(\pixelfeed/N166 ) );
  GTECH_AND2 \pixelfeed/C280  ( .A(\pixelfeed/N161 ), .B(\pixelfeed/N162 ), 
        .Z(\pixelfeed/N165 ) );
  \**SEQGEN**  \pixelfeed/ignore_reg  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N157 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\pixelfeed/ignore ), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N156 ) );
  \**SEQGEN**  \pixelfeed/state_reg_0_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N152 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\pixelfeed/state[0] ), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N226 ) );
  \**SEQGEN**  \pixelfeed/state_reg_1_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N153 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\pixelfeed/state[1] ), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N226 ) );
  \**SEQGEN**  \pixelfeed/state_reg_2_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N154 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\pixelfeed/state[2] ), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N226 ) );
  \**SEQGEN**  \pixelfeed/state_reg_3_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N155 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\pixelfeed/state[3] ), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N226 ) );
  \**SEQGEN**  \pixelfeed/dcb_index_reg_0_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N149 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(dcb_adr[3]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \pixelfeed/dcb_index_reg_1_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N150 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(dcb_adr[4]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_0_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N118 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[0]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_1_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N119 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[1]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_2_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N120 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[2]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_3_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N121 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[3]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_4_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N122 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[4]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_5_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N123 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[5]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_6_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N124 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[6]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_7_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N125 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[7]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_8_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N126 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[8]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_9_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N127 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[9]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_10_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N128 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[10]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_11_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N129 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[11]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_12_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N130 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[12]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_13_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N131 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[13]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_14_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N132 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[14]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_15_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N133 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[15]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_16_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N134 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[16]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_17_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N135 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[17]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_18_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N136 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[18]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_19_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N137 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[19]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_20_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N138 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[20]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_21_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N139 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[21]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_22_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N140 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[22]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_23_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N141 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[23]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_24_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N142 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[24]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/fml_adr_reg_25_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N143 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(fml_adr[25]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N117 ) );
  \**SEQGEN**  \pixelfeed/sof_reg  ( .clear(1'b0), .preset(1'b0), .next_state(
        \pixelfeed/N60 ), .clocked_on(sys_clk), .data_in(1'b0), .enable(1'b0), 
        .Q(\pixelfeed/sof ), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(\pixelfeed/N41 ) );
  \**SEQGEN**  \pixelfeed/bcounter_reg_0_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N42 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\pixelfeed/bcounter[0] ), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N41 ) );
  \**SEQGEN**  \pixelfeed/bcounter_reg_1_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N43 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\pixelfeed/bcounter[1] ), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N41 ) );
  \**SEQGEN**  \pixelfeed/bcounter_reg_2_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N44 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\pixelfeed/bcounter[2] ), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N41 ) );
  \**SEQGEN**  \pixelfeed/bcounter_reg_3_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N45 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\pixelfeed/bcounter[3] ), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N41 ) );
  \**SEQGEN**  \pixelfeed/bcounter_reg_4_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N46 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\pixelfeed/bcounter[4] ), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N41 ) );
  \**SEQGEN**  \pixelfeed/bcounter_reg_5_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N47 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\pixelfeed/bcounter[5] ), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N41 ) );
  \**SEQGEN**  \pixelfeed/bcounter_reg_6_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N48 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\pixelfeed/bcounter[6] ), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N41 ) );
  \**SEQGEN**  \pixelfeed/bcounter_reg_7_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N49 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\pixelfeed/bcounter[7] ), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N41 ) );
  \**SEQGEN**  \pixelfeed/bcounter_reg_8_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N50 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\pixelfeed/bcounter[8] ), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N41 ) );
  \**SEQGEN**  \pixelfeed/bcounter_reg_9_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N51 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\pixelfeed/bcounter[9] ), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N41 ) );
  \**SEQGEN**  \pixelfeed/bcounter_reg_10_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N52 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\pixelfeed/bcounter[10] ), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N41 ) );
  \**SEQGEN**  \pixelfeed/bcounter_reg_11_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N53 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\pixelfeed/bcounter[11] ), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N41 ) );
  \**SEQGEN**  \pixelfeed/bcounter_reg_12_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N54 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\pixelfeed/bcounter[12] ), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N41 ) );
  \**SEQGEN**  \pixelfeed/bcounter_reg_13_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N55 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\pixelfeed/bcounter[13] ), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N41 ) );
  \**SEQGEN**  \pixelfeed/bcounter_reg_14_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N56 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\pixelfeed/bcounter[14] ), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N41 ) );
  \**SEQGEN**  \pixelfeed/bcounter_reg_15_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N57 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\pixelfeed/bcounter[15] ), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N41 ) );
  \**SEQGEN**  \pixelfeed/bcounter_reg_16_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N58 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\pixelfeed/bcounter[16] ), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N41 ) );
  \**SEQGEN**  \pixelfeed/bcounter_reg_17_  ( .clear(1'b0), .preset(1'b0), 
        .next_state(\pixelfeed/N59 ), .clocked_on(sys_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(\pixelfeed/bcounter[17] ), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/N41 ) );
  EQ_UNS_OP \pixelfeed/eq_80  ( .A({\pixelfeed/bcounter[17] , 
        \pixelfeed/bcounter[16] , \pixelfeed/bcounter[15] , 
        \pixelfeed/bcounter[14] , \pixelfeed/bcounter[13] , 
        \pixelfeed/bcounter[12] , \pixelfeed/bcounter[11] , 
        \pixelfeed/bcounter[10] , \pixelfeed/bcounter[9] , 
        \pixelfeed/bcounter[8] , \pixelfeed/bcounter[7] , 
        \pixelfeed/bcounter[6] , \pixelfeed/bcounter[5] , 
        \pixelfeed/bcounter[4] , \pixelfeed/bcounter[3] , 
        \pixelfeed/bcounter[2] , \pixelfeed/bcounter[1] , 
        \pixelfeed/bcounter[0] }), .B(nbursts), .Z(\pixelfeed/N38 ) );
  GTECH_NOT \pixelfeed/fifo64to16/I_12  ( .A(\pixelfeed/fifo64to16/N81 ), .Z(
        pixel_valid) );
  GTECH_AND2 \pixelfeed/fifo64to16/C1744  ( .A(\pixelfeed/fifo64to16/N25 ), 
        .B(pixel_ack), .Z() );
  GTECH_NOT \pixelfeed/fifo64to16/I_11  ( .A(pixel_ack), .Z(
        \pixelfeed/fifo64to16/N43 ) );
  GTECH_AND2 \pixelfeed/fifo64to16/C1739  ( .A(\pixelfeed/fifo64to16/N26 ), 
        .B(\pixelfeed/fifo64to16/level[0] ), .Z(\pixelfeed/fifo64to16/N95 ) );
  GTECH_AND2 \pixelfeed/fifo64to16/C1738  ( .A(\pixelfeed/fifo_stb ), .B(
        \pixelfeed/fifo64to16/N29 ), .Z(\pixelfeed/fifo64to16/N94 ) );
  GTECH_OR2 \pixelfeed/fifo64to16/C1737  ( .A(\pixelfeed/fifo64to16/N94 ), .B(
        \pixelfeed/fifo64to16/N95 ), .Z(\pixelfeed/fifo64to16/N42 ) );
  GTECH_AND2 \pixelfeed/fifo64to16/C1735  ( .A(\pixelfeed/fifo64to16/N26 ), 
        .B(\pixelfeed/fifo64to16/level[1] ), .Z(\pixelfeed/fifo64to16/N93 ) );
  GTECH_AND2 \pixelfeed/fifo64to16/C1734  ( .A(\pixelfeed/fifo_stb ), .B(
        \pixelfeed/fifo64to16/N30 ), .Z(\pixelfeed/fifo64to16/N92 ) );
  GTECH_OR2 \pixelfeed/fifo64to16/C1733  ( .A(\pixelfeed/fifo64to16/N92 ), .B(
        \pixelfeed/fifo64to16/N93 ), .Z(\pixelfeed/fifo64to16/N41 ) );
  GTECH_AND2 \pixelfeed/fifo64to16/C1731  ( .A(\pixelfeed/fifo64to16/N26 ), 
        .B(\pixelfeed/fifo64to16/level[2] ), .Z(\pixelfeed/fifo64to16/N91 ) );
  GTECH_AND2 \pixelfeed/fifo64to16/C1730  ( .A(\pixelfeed/fifo_stb ), .B(
        \pixelfeed/fifo64to16/N31 ), .Z(\pixelfeed/fifo64to16/N90 ) );
  GTECH_OR2 \pixelfeed/fifo64to16/C1729  ( .A(\pixelfeed/fifo64to16/N90 ), .B(
        \pixelfeed/fifo64to16/N91 ), .Z(\pixelfeed/fifo64to16/N40 ) );
  GTECH_AND2 \pixelfeed/fifo64to16/C1727  ( .A(\pixelfeed/fifo64to16/N26 ), 
        .B(\pixelfeed/fifo64to16/level[3] ), .Z(\pixelfeed/fifo64to16/N89 ) );
  GTECH_AND2 \pixelfeed/fifo64to16/C1726  ( .A(\pixelfeed/fifo_stb ), .B(
        \pixelfeed/fifo64to16/N32 ), .Z(\pixelfeed/fifo64to16/N88 ) );
  GTECH_OR2 \pixelfeed/fifo64to16/C1725  ( .A(\pixelfeed/fifo64to16/N88 ), .B(
        \pixelfeed/fifo64to16/N89 ), .Z(\pixelfeed/fifo64to16/N39 ) );
  GTECH_AND2 \pixelfeed/fifo64to16/C1723  ( .A(\pixelfeed/fifo64to16/N26 ), 
        .B(\pixelfeed/fifo64to16/level[4] ), .Z(\pixelfeed/fifo64to16/N87 ) );
  GTECH_AND2 \pixelfeed/fifo64to16/C1722  ( .A(\pixelfeed/fifo_stb ), .B(
        \pixelfeed/fifo64to16/N33 ), .Z(\pixelfeed/fifo64to16/N86 ) );
  GTECH_OR2 \pixelfeed/fifo64to16/C1721  ( .A(\pixelfeed/fifo64to16/N86 ), .B(
        \pixelfeed/fifo64to16/N87 ), .Z(\pixelfeed/fifo64to16/N38 ) );
  GTECH_AND2 \pixelfeed/fifo64to16/C1716  ( .A(\pixelfeed/fifo64to16/N25 ), 
        .B(\pixelfeed/fifo_stb ), .Z() );
  GTECH_NOT \pixelfeed/fifo64to16/I_10  ( .A(\pixelfeed/fifo_stb ), .Z(
        \pixelfeed/fifo64to16/N26 ) );
  GTECH_BUF \pixelfeed/fifo64to16/B_12  ( .A(\pixelfeed/fifo64to16/N24 ), .Z(
        \pixelfeed/fifo64to16/N25 ) );
  GTECH_NOT \pixelfeed/fifo64to16/I_9  ( .A(vga_rst), .Z(
        \pixelfeed/fifo64to16/N24 ) );
  GTECH_NOT \pixelfeed/fifo64to16/I_8  ( .A(\pixelfeed/fifo64to16/N21 ), .Z(
        \pixelfeed/fifo64to16/N22 ) );
  GTECH_NOT \pixelfeed/fifo64to16/I_7  ( .A(\pixelfeed/fifo64to16/N19 ), .Z(
        \pixelfeed/fifo64to16/N20 ) );
  GTECH_NOT \pixelfeed/fifo64to16/I_6  ( .A(\pixelfeed/fifo64to16/consume[0] ), 
        .Z(\pixelfeed/fifo64to16/N17 ) );
  GTECH_NOT \pixelfeed/fifo64to16/I_5  ( .A(\pixelfeed/fifo64to16/consume[1] ), 
        .Z(\pixelfeed/fifo64to16/N16 ) );
  GTECH_BUF \pixelfeed/fifo64to16/B_11  ( .A(\pixelfeed/fifo64to16/consume[3] ), .Z(\pixelfeed/fifo64to16/N15 ) );
  GTECH_BUF \pixelfeed/fifo64to16/B_10  ( .A(\pixelfeed/fifo64to16/consume[2] ), .Z(\pixelfeed/fifo64to16/N14 ) );
  MUX_OP \pixelfeed/fifo64to16/C1696  ( .D0({
        \pixelfeed/fifo64to16/storage  [192], 
        \pixelfeed/fifo64to16/storage  [193], 
        \pixelfeed/fifo64to16/storage  [194], 
        \pixelfeed/fifo64to16/storage  [195], 
        \pixelfeed/fifo64to16/storage  [196], 
        \pixelfeed/fifo64to16/storage  [197], 
        \pixelfeed/fifo64to16/storage  [198], 
        \pixelfeed/fifo64to16/storage  [199], 
        \pixelfeed/fifo64to16/storage  [200], 
        \pixelfeed/fifo64to16/storage  [201], 
        \pixelfeed/fifo64to16/storage  [202], 
        \pixelfeed/fifo64to16/storage  [203], 
        \pixelfeed/fifo64to16/storage  [204], 
        \pixelfeed/fifo64to16/storage  [205], 
        \pixelfeed/fifo64to16/storage  [206], 
        \pixelfeed/fifo64to16/storage  [207], 
        \pixelfeed/fifo64to16/storage  [208], 
        \pixelfeed/fifo64to16/storage  [209], 
        \pixelfeed/fifo64to16/storage  [210], 
        \pixelfeed/fifo64to16/storage  [211], 
        \pixelfeed/fifo64to16/storage  [212], 
        \pixelfeed/fifo64to16/storage  [213], 
        \pixelfeed/fifo64to16/storage  [214], 
        \pixelfeed/fifo64to16/storage  [215], 
        \pixelfeed/fifo64to16/storage  [216], 
        \pixelfeed/fifo64to16/storage  [217], 
        \pixelfeed/fifo64to16/storage  [218], 
        \pixelfeed/fifo64to16/storage  [219], 
        \pixelfeed/fifo64to16/storage  [220], 
        \pixelfeed/fifo64to16/storage  [221], 
        \pixelfeed/fifo64to16/storage  [222], 
        \pixelfeed/fifo64to16/storage  [223], 
        \pixelfeed/fifo64to16/storage  [224], 
        \pixelfeed/fifo64to16/storage  [225], 
        \pixelfeed/fifo64to16/storage  [226], 
        \pixelfeed/fifo64to16/storage  [227], 
        \pixelfeed/fifo64to16/storage  [228], 
        \pixelfeed/fifo64to16/storage  [229], 
        \pixelfeed/fifo64to16/storage  [230], 
        \pixelfeed/fifo64to16/storage  [231], 
        \pixelfeed/fifo64to16/storage  [232], 
        \pixelfeed/fifo64to16/storage  [233], 
        \pixelfeed/fifo64to16/storage  [234], 
        \pixelfeed/fifo64to16/storage  [235], 
        \pixelfeed/fifo64to16/storage  [236], 
        \pixelfeed/fifo64to16/storage  [237], 
        \pixelfeed/fifo64to16/storage  [238], 
        \pixelfeed/fifo64to16/storage  [239], 
        \pixelfeed/fifo64to16/storage  [240], 
        \pixelfeed/fifo64to16/storage  [241], 
        \pixelfeed/fifo64to16/storage  [242], 
        \pixelfeed/fifo64to16/storage  [243], 
        \pixelfeed/fifo64to16/storage  [244], 
        \pixelfeed/fifo64to16/storage  [245], 
        \pixelfeed/fifo64to16/storage  [246], 
        \pixelfeed/fifo64to16/storage  [247], 
        \pixelfeed/fifo64to16/storage  [248], 
        \pixelfeed/fifo64to16/storage  [249], 
        \pixelfeed/fifo64to16/storage  [250], 
        \pixelfeed/fifo64to16/storage  [251], 
        \pixelfeed/fifo64to16/storage  [252], 
        \pixelfeed/fifo64to16/storage  [253], 
        \pixelfeed/fifo64to16/storage  [254], 
        \pixelfeed/fifo64to16/storage  [255]}), .D1({
        \pixelfeed/fifo64to16/storage  [128], 
        \pixelfeed/fifo64to16/storage  [129], 
        \pixelfeed/fifo64to16/storage  [130], 
        \pixelfeed/fifo64to16/storage  [131], 
        \pixelfeed/fifo64to16/storage  [132], 
        \pixelfeed/fifo64to16/storage  [133], 
        \pixelfeed/fifo64to16/storage  [134], 
        \pixelfeed/fifo64to16/storage  [135], 
        \pixelfeed/fifo64to16/storage  [136], 
        \pixelfeed/fifo64to16/storage  [137], 
        \pixelfeed/fifo64to16/storage  [138], 
        \pixelfeed/fifo64to16/storage  [139], 
        \pixelfeed/fifo64to16/storage  [140], 
        \pixelfeed/fifo64to16/storage  [141], 
        \pixelfeed/fifo64to16/storage  [142], 
        \pixelfeed/fifo64to16/storage  [143], 
        \pixelfeed/fifo64to16/storage  [144], 
        \pixelfeed/fifo64to16/storage  [145], 
        \pixelfeed/fifo64to16/storage  [146], 
        \pixelfeed/fifo64to16/storage  [147], 
        \pixelfeed/fifo64to16/storage  [148], 
        \pixelfeed/fifo64to16/storage  [149], 
        \pixelfeed/fifo64to16/storage  [150], 
        \pixelfeed/fifo64to16/storage  [151], 
        \pixelfeed/fifo64to16/storage  [152], 
        \pixelfeed/fifo64to16/storage  [153], 
        \pixelfeed/fifo64to16/storage  [154], 
        \pixelfeed/fifo64to16/storage  [155], 
        \pixelfeed/fifo64to16/storage  [156], 
        \pixelfeed/fifo64to16/storage  [157], 
        \pixelfeed/fifo64to16/storage  [158], 
        \pixelfeed/fifo64to16/storage  [159], 
        \pixelfeed/fifo64to16/storage  [160], 
        \pixelfeed/fifo64to16/storage  [161], 
        \pixelfeed/fifo64to16/storage  [162], 
        \pixelfeed/fifo64to16/storage  [163], 
        \pixelfeed/fifo64to16/storage  [164], 
        \pixelfeed/fifo64to16/storage  [165], 
        \pixelfeed/fifo64to16/storage  [166], 
        \pixelfeed/fifo64to16/storage  [167], 
        \pixelfeed/fifo64to16/storage  [168], 
        \pixelfeed/fifo64to16/storage  [169], 
        \pixelfeed/fifo64to16/storage  [170], 
        \pixelfeed/fifo64to16/storage  [171], 
        \pixelfeed/fifo64to16/storage  [172], 
        \pixelfeed/fifo64to16/storage  [173], 
        \pixelfeed/fifo64to16/storage  [174], 
        \pixelfeed/fifo64to16/storage  [175], 
        \pixelfeed/fifo64to16/storage  [176], 
        \pixelfeed/fifo64to16/storage  [177], 
        \pixelfeed/fifo64to16/storage  [178], 
        \pixelfeed/fifo64to16/storage  [179], 
        \pixelfeed/fifo64to16/storage  [180], 
        \pixelfeed/fifo64to16/storage  [181], 
        \pixelfeed/fifo64to16/storage  [182], 
        \pixelfeed/fifo64to16/storage  [183], 
        \pixelfeed/fifo64to16/storage  [184], 
        \pixelfeed/fifo64to16/storage  [185], 
        \pixelfeed/fifo64to16/storage  [186], 
        \pixelfeed/fifo64to16/storage  [187], 
        \pixelfeed/fifo64to16/storage  [188], 
        \pixelfeed/fifo64to16/storage  [189], 
        \pixelfeed/fifo64to16/storage  [190], 
        \pixelfeed/fifo64to16/storage  [191]}), .D2({
        \pixelfeed/fifo64to16/storage  [64], 
        \pixelfeed/fifo64to16/storage  [65], 
        \pixelfeed/fifo64to16/storage  [66], 
        \pixelfeed/fifo64to16/storage  [67], 
        \pixelfeed/fifo64to16/storage  [68], 
        \pixelfeed/fifo64to16/storage  [69], 
        \pixelfeed/fifo64to16/storage  [70], 
        \pixelfeed/fifo64to16/storage  [71], 
        \pixelfeed/fifo64to16/storage  [72], 
        \pixelfeed/fifo64to16/storage  [73], 
        \pixelfeed/fifo64to16/storage  [74], 
        \pixelfeed/fifo64to16/storage  [75], 
        \pixelfeed/fifo64to16/storage  [76], 
        \pixelfeed/fifo64to16/storage  [77], 
        \pixelfeed/fifo64to16/storage  [78], 
        \pixelfeed/fifo64to16/storage  [79], 
        \pixelfeed/fifo64to16/storage  [80], 
        \pixelfeed/fifo64to16/storage  [81], 
        \pixelfeed/fifo64to16/storage  [82], 
        \pixelfeed/fifo64to16/storage  [83], 
        \pixelfeed/fifo64to16/storage  [84], 
        \pixelfeed/fifo64to16/storage  [85], 
        \pixelfeed/fifo64to16/storage  [86], 
        \pixelfeed/fifo64to16/storage  [87], 
        \pixelfeed/fifo64to16/storage  [88], 
        \pixelfeed/fifo64to16/storage  [89], 
        \pixelfeed/fifo64to16/storage  [90], 
        \pixelfeed/fifo64to16/storage  [91], 
        \pixelfeed/fifo64to16/storage  [92], 
        \pixelfeed/fifo64to16/storage  [93], 
        \pixelfeed/fifo64to16/storage  [94], 
        \pixelfeed/fifo64to16/storage  [95], 
        \pixelfeed/fifo64to16/storage  [96], 
        \pixelfeed/fifo64to16/storage  [97], 
        \pixelfeed/fifo64to16/storage  [98], 
        \pixelfeed/fifo64to16/storage  [99], 
        \pixelfeed/fifo64to16/storage  [100], 
        \pixelfeed/fifo64to16/storage  [101], 
        \pixelfeed/fifo64to16/storage  [102], 
        \pixelfeed/fifo64to16/storage  [103], 
        \pixelfeed/fifo64to16/storage  [104], 
        \pixelfeed/fifo64to16/storage  [105], 
        \pixelfeed/fifo64to16/storage  [106], 
        \pixelfeed/fifo64to16/storage  [107], 
        \pixelfeed/fifo64to16/storage  [108], 
        \pixelfeed/fifo64to16/storage  [109], 
        \pixelfeed/fifo64to16/storage  [110], 
        \pixelfeed/fifo64to16/storage  [111], 
        \pixelfeed/fifo64to16/storage  [112], 
        \pixelfeed/fifo64to16/storage  [113], 
        \pixelfeed/fifo64to16/storage  [114], 
        \pixelfeed/fifo64to16/storage  [115], 
        \pixelfeed/fifo64to16/storage  [116], 
        \pixelfeed/fifo64to16/storage  [117], 
        \pixelfeed/fifo64to16/storage  [118], 
        \pixelfeed/fifo64to16/storage  [119], 
        \pixelfeed/fifo64to16/storage  [120], 
        \pixelfeed/fifo64to16/storage  [121], 
        \pixelfeed/fifo64to16/storage  [122], 
        \pixelfeed/fifo64to16/storage  [123], 
        \pixelfeed/fifo64to16/storage  [124], 
        \pixelfeed/fifo64to16/storage  [125], 
        \pixelfeed/fifo64to16/storage  [126], 
        \pixelfeed/fifo64to16/storage  [127]}), .D3({
        \pixelfeed/fifo64to16/storage  [0], \pixelfeed/fifo64to16/storage  [1], 
        \pixelfeed/fifo64to16/storage  [2], \pixelfeed/fifo64to16/storage  [3], 
        \pixelfeed/fifo64to16/storage  [4], \pixelfeed/fifo64to16/storage  [5], 
        \pixelfeed/fifo64to16/storage  [6], \pixelfeed/fifo64to16/storage  [7], 
        \pixelfeed/fifo64to16/storage  [8], \pixelfeed/fifo64to16/storage  [9], 
        \pixelfeed/fifo64to16/storage  [10], 
        \pixelfeed/fifo64to16/storage  [11], 
        \pixelfeed/fifo64to16/storage  [12], 
        \pixelfeed/fifo64to16/storage  [13], 
        \pixelfeed/fifo64to16/storage  [14], 
        \pixelfeed/fifo64to16/storage  [15], 
        \pixelfeed/fifo64to16/storage  [16], 
        \pixelfeed/fifo64to16/storage  [17], 
        \pixelfeed/fifo64to16/storage  [18], 
        \pixelfeed/fifo64to16/storage  [19], 
        \pixelfeed/fifo64to16/storage  [20], 
        \pixelfeed/fifo64to16/storage  [21], 
        \pixelfeed/fifo64to16/storage  [22], 
        \pixelfeed/fifo64to16/storage  [23], 
        \pixelfeed/fifo64to16/storage  [24], 
        \pixelfeed/fifo64to16/storage  [25], 
        \pixelfeed/fifo64to16/storage  [26], 
        \pixelfeed/fifo64to16/storage  [27], 
        \pixelfeed/fifo64to16/storage  [28], 
        \pixelfeed/fifo64to16/storage  [29], 
        \pixelfeed/fifo64to16/storage  [30], 
        \pixelfeed/fifo64to16/storage  [31], 
        \pixelfeed/fifo64to16/storage  [32], 
        \pixelfeed/fifo64to16/storage  [33], 
        \pixelfeed/fifo64to16/storage  [34], 
        \pixelfeed/fifo64to16/storage  [35], 
        \pixelfeed/fifo64to16/storage  [36], 
        \pixelfeed/fifo64to16/storage  [37], 
        \pixelfeed/fifo64to16/storage  [38], 
        \pixelfeed/fifo64to16/storage  [39], 
        \pixelfeed/fifo64to16/storage  [40], 
        \pixelfeed/fifo64to16/storage  [41], 
        \pixelfeed/fifo64to16/storage  [42], 
        \pixelfeed/fifo64to16/storage  [43], 
        \pixelfeed/fifo64to16/storage  [44], 
        \pixelfeed/fifo64to16/storage  [45], 
        \pixelfeed/fifo64to16/storage  [46], 
        \pixelfeed/fifo64to16/storage  [47], 
        \pixelfeed/fifo64to16/storage  [48], 
        \pixelfeed/fifo64to16/storage  [49], 
        \pixelfeed/fifo64to16/storage  [50], 
        \pixelfeed/fifo64to16/storage  [51], 
        \pixelfeed/fifo64to16/storage  [52], 
        \pixelfeed/fifo64to16/storage  [53], 
        \pixelfeed/fifo64to16/storage  [54], 
        \pixelfeed/fifo64to16/storage  [55], 
        \pixelfeed/fifo64to16/storage  [56], 
        \pixelfeed/fifo64to16/storage  [57], 
        \pixelfeed/fifo64to16/storage  [58], 
        \pixelfeed/fifo64to16/storage  [59], 
        \pixelfeed/fifo64to16/storage  [60], 
        \pixelfeed/fifo64to16/storage  [61], 
        \pixelfeed/fifo64to16/storage  [62], 
        \pixelfeed/fifo64to16/storage  [63]}), .S0(\pixelfeed/fifo64to16/N14 ), 
        .S1(\pixelfeed/fifo64to16/N15 ), .Z({\pixelfeed/fifo64to16/do64  [0], 
        \pixelfeed/fifo64to16/do64  [1], \pixelfeed/fifo64to16/do64  [2], 
        \pixelfeed/fifo64to16/do64  [3], \pixelfeed/fifo64to16/do64  [4], 
        \pixelfeed/fifo64to16/do64  [5], \pixelfeed/fifo64to16/do64  [6], 
        \pixelfeed/fifo64to16/do64  [7], \pixelfeed/fifo64to16/do64  [8], 
        \pixelfeed/fifo64to16/do64  [9], \pixelfeed/fifo64to16/do64  [10], 
        \pixelfeed/fifo64to16/do64  [11], \pixelfeed/fifo64to16/do64  [12], 
        \pixelfeed/fifo64to16/do64  [13], \pixelfeed/fifo64to16/do64  [14], 
        \pixelfeed/fifo64to16/do64  [15], \pixelfeed/fifo64to16/do64  [16], 
        \pixelfeed/fifo64to16/do64  [17], \pixelfeed/fifo64to16/do64  [18], 
        \pixelfeed/fifo64to16/do64  [19], \pixelfeed/fifo64to16/do64  [20], 
        \pixelfeed/fifo64to16/do64  [21], \pixelfeed/fifo64to16/do64  [22], 
        \pixelfeed/fifo64to16/do64  [23], \pixelfeed/fifo64to16/do64  [24], 
        \pixelfeed/fifo64to16/do64  [25], \pixelfeed/fifo64to16/do64  [26], 
        \pixelfeed/fifo64to16/do64  [27], \pixelfeed/fifo64to16/do64  [28], 
        \pixelfeed/fifo64to16/do64  [29], \pixelfeed/fifo64to16/do64  [30], 
        \pixelfeed/fifo64to16/do64  [31], \pixelfeed/fifo64to16/do64  [32], 
        \pixelfeed/fifo64to16/do64  [33], \pixelfeed/fifo64to16/do64  [34], 
        \pixelfeed/fifo64to16/do64  [35], \pixelfeed/fifo64to16/do64  [36], 
        \pixelfeed/fifo64to16/do64  [37], \pixelfeed/fifo64to16/do64  [38], 
        \pixelfeed/fifo64to16/do64  [39], \pixelfeed/fifo64to16/do64  [40], 
        \pixelfeed/fifo64to16/do64  [41], \pixelfeed/fifo64to16/do64  [42], 
        \pixelfeed/fifo64to16/do64  [43], \pixelfeed/fifo64to16/do64  [44], 
        \pixelfeed/fifo64to16/do64  [45], \pixelfeed/fifo64to16/do64  [46], 
        \pixelfeed/fifo64to16/do64  [47], \pixelfeed/fifo64to16/do64  [48], 
        \pixelfeed/fifo64to16/do64  [49], \pixelfeed/fifo64to16/do64  [50], 
        \pixelfeed/fifo64to16/do64  [51], \pixelfeed/fifo64to16/do64  [52], 
        \pixelfeed/fifo64to16/do64  [53], \pixelfeed/fifo64to16/do64  [54], 
        \pixelfeed/fifo64to16/do64  [55], \pixelfeed/fifo64to16/do64  [56], 
        \pixelfeed/fifo64to16/do64  [57], \pixelfeed/fifo64to16/do64  [58], 
        \pixelfeed/fifo64to16/do64  [59], \pixelfeed/fifo64to16/do64  [60], 
        \pixelfeed/fifo64to16/do64  [61], \pixelfeed/fifo64to16/do64  [62], 
        \pixelfeed/fifo64to16/do64  [63]}) );
  SELECT_OP \pixelfeed/fifo64to16/C1695  ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2({\pixelfeed/fifo64to16/N37 , \pixelfeed/fifo64to16/N36 , 
        \pixelfeed/fifo64to16/N35 , \pixelfeed/fifo64to16/N34 }), .CONTROL1(
        \pixelfeed/fifo64to16/N12 ), .CONTROL2(\pixelfeed/fifo64to16/N13 ), 
        .Z({\pixelfeed/fifo64to16/N76 , \pixelfeed/fifo64to16/N75 , 
        \pixelfeed/fifo64to16/N74 , \pixelfeed/fifo64to16/N73 }) );
  SELECT_OP \pixelfeed/fifo64to16/C1694  ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .DATA2({\pixelfeed/fifo64to16/N58 , \pixelfeed/fifo64to16/N57 , 
        \pixelfeed/fifo64to16/N56 , \pixelfeed/fifo64to16/N55 , 
        \pixelfeed/fifo64to16/N54 }), .CONTROL1(\pixelfeed/fifo64to16/N12 ), 
        .CONTROL2(\pixelfeed/fifo64to16/N13 ), .Z({\pixelfeed/fifo64to16/N72 , 
        \pixelfeed/fifo64to16/N71 , \pixelfeed/fifo64to16/N70 , 
        \pixelfeed/fifo64to16/N69 , \pixelfeed/fifo64to16/N68 }) );
  SELECT_OP \pixelfeed/fifo64to16/C1693  ( .DATA1(1'b1), .DATA2(
        \pixelfeed/fifo64to16/N53 ), .CONTROL1(\pixelfeed/fifo64to16/N12 ), 
        .CONTROL2(\pixelfeed/fifo64to16/N13 ), .Z(\pixelfeed/fifo64to16/N67 )
         );
  SELECT_OP \pixelfeed/fifo64to16/C1692  ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2({\pixelfeed/fifo64to16/N47 , \pixelfeed/fifo64to16/N46 , 
        \pixelfeed/fifo64to16/N45 , \pixelfeed/fifo64to16/N44 }), .CONTROL1(
        \pixelfeed/fifo64to16/N12 ), .CONTROL2(\pixelfeed/fifo64to16/N13 ), 
        .Z({\pixelfeed/fifo64to16/N66 , \pixelfeed/fifo64to16/N65 , 
        \pixelfeed/fifo64to16/N64 , \pixelfeed/fifo64to16/N63 }) );
  SELECT_OP \pixelfeed/fifo64to16/C1691  ( .DATA1(1'b1), .DATA2(pixel_ack), 
        .CONTROL1(\pixelfeed/fifo64to16/N12 ), .CONTROL2(
        \pixelfeed/fifo64to16/N13 ), .Z(\pixelfeed/fifo64to16/N62 ) );
  SELECT_OP \pixelfeed/fifo64to16/C1690  ( .DATA1({1'b0, 1'b0}), .DATA2({
        \pixelfeed/fifo64to16/N28 , \pixelfeed/fifo64to16/N27 }), .CONTROL1(
        \pixelfeed/fifo64to16/N12 ), .CONTROL2(\pixelfeed/fifo64to16/N13 ), 
        .Z({\pixelfeed/fifo64to16/N61 , \pixelfeed/fifo64to16/N60 }) );
  GTECH_BUF \pixelfeed/fifo64to16/B_9  ( .A(\pixelfeed/fifo64to16/N24 ), .Z(
        \pixelfeed/fifo64to16/N13 ) );
  GTECH_BUF \pixelfeed/fifo64to16/B_8  ( .A(vga_rst), .Z(
        \pixelfeed/fifo64to16/N12 ) );
  SELECT_OP \pixelfeed/fifo64to16/C1689  ( .DATA1(1'b1), .DATA2(
        \pixelfeed/fifo_stb ), .CONTROL1(\pixelfeed/fifo64to16/N12 ), 
        .CONTROL2(\pixelfeed/fifo64to16/N13 ), .Z(\pixelfeed/fifo64to16/N59 )
         );
  SELECT_OP \pixelfeed/fifo64to16/C1688  ( .DATA1({\pixelfeed/fifo64to16/N52 , 
        \pixelfeed/fifo64to16/N51 , \pixelfeed/fifo64to16/N50 , 
        \pixelfeed/fifo64to16/N49 , \pixelfeed/fifo64to16/N48 }), .DATA2({
        \pixelfeed/fifo64to16/N33 , \pixelfeed/fifo64to16/N32 , 
        \pixelfeed/fifo64to16/N31 , \pixelfeed/fifo64to16/N30 , 
        \pixelfeed/fifo64to16/N29 }), .CONTROL1(\pixelfeed/fifo64to16/N10 ), 
        .CONTROL2(\pixelfeed/fifo64to16/N11 ), .Z({\pixelfeed/fifo64to16/N58 , 
        \pixelfeed/fifo64to16/N57 , \pixelfeed/fifo64to16/N56 , 
        \pixelfeed/fifo64to16/N55 , \pixelfeed/fifo64to16/N54 }) );
  GTECH_BUF \pixelfeed/fifo64to16/B_7  ( .A(\pixelfeed/fifo64to16/N43 ), .Z(
        \pixelfeed/fifo64to16/N11 ) );
  GTECH_BUF \pixelfeed/fifo64to16/B_6  ( .A(pixel_ack), .Z(
        \pixelfeed/fifo64to16/N10 ) );
  SELECT_OP \pixelfeed/fifo64to16/C1687  ( .DATA1(1'b1), .DATA2(
        \pixelfeed/fifo_stb ), .CONTROL1(\pixelfeed/fifo64to16/N10 ), 
        .CONTROL2(\pixelfeed/fifo64to16/N11 ), .Z(\pixelfeed/fifo64to16/N53 )
         );
  GTECH_BUF \pixelfeed/fifo64to16/B_5  ( .A(\pixelfeed/fifo64to16/N26 ), .Z(
        \pixelfeed/fifo64to16/N9 ) );
  GTECH_BUF \pixelfeed/fifo64to16/B_4  ( .A(\pixelfeed/fifo_stb ), .Z(
        \pixelfeed/fifo64to16/N8 ) );
  SELECT_OP \pixelfeed/fifo64to16/C1686  ( .DATA1({\pixelfeed/fifo64to16/N85 , 
        \pixelfeed/fifo64to16/N84 , \pixelfeed/fifo64to16/N83 , 
        \pixelfeed/fifo64to16/N82 }), .DATA2({1'b0, 1'b0, 1'b0, 1'b0}), 
        .CONTROL1(\pixelfeed/fifo64to16/N8 ), .CONTROL2(
        \pixelfeed/fifo64to16/N9 ), .Z({\pixelfeed/fifo64to16/N37 , 
        \pixelfeed/fifo64to16/N36 , \pixelfeed/fifo64to16/N35 , 
        \pixelfeed/fifo64to16/N34 }) );
  GTECH_BUF \pixelfeed/fifo64to16/B_3  ( .A(\pixelfeed/fifo64to16/N23 ), .Z(
        \pixelfeed/fifo64to16/N7 ) );
  GTECH_BUF \pixelfeed/fifo64to16/B_2  ( .A(\pixelfeed/fifo64to16/N22 ), .Z(
        \pixelfeed/fifo64to16/N6 ) );
  GTECH_BUF \pixelfeed/fifo64to16/B_1  ( .A(\pixelfeed/fifo64to16/N20 ), .Z(
        \pixelfeed/fifo64to16/N5 ) );
  GTECH_BUF \pixelfeed/fifo64to16/B_0  ( .A(\pixelfeed/fifo64to16/N18 ), .Z(
        \pixelfeed/fifo64to16/N4 ) );
  SELECT_OP \pixelfeed/fifo64to16/C1685  ( .DATA1(
        \pixelfeed/fifo64to16/do64 [63:48]), .DATA2(
        \pixelfeed/fifo64to16/do64 [47:32]), .DATA3(
        \pixelfeed/fifo64to16/do64 [31:16]), .DATA4(
        \pixelfeed/fifo64to16/do64 [15:0]), .CONTROL1(
        \pixelfeed/fifo64to16/N4 ), .CONTROL2(\pixelfeed/fifo64to16/N5 ), 
        .CONTROL3(\pixelfeed/fifo64to16/N6 ), .CONTROL4(
        \pixelfeed/fifo64to16/N7 ), .Z(pixel_fb) );
  GTECH_NOT \pixelfeed/fifo64to16/I_4  ( .A(\pixelfeed/fifo64to16/produce[1] ), 
        .Z(\pixelfeed/fifo64to16/N3 ) );
  GTECH_NOT \pixelfeed/fifo64to16/I_3  ( .A(\pixelfeed/fifo64to16/produce[0] ), 
        .Z(\pixelfeed/fifo64to16/N2 ) );
  GTECH_AND2 \pixelfeed/fifo64to16/C1684  ( .A(\pixelfeed/fifo64to16/N2 ), .B(
        \pixelfeed/fifo64to16/N3 ), .Z(\pixelfeed/fifo64to16/N85 ) );
  GTECH_NOT \pixelfeed/fifo64to16/I_2  ( .A(\pixelfeed/fifo64to16/produce[1] ), 
        .Z(\pixelfeed/fifo64to16/N1 ) );
  GTECH_AND2 \pixelfeed/fifo64to16/C1683  ( .A(
        \pixelfeed/fifo64to16/produce[0] ), .B(\pixelfeed/fifo64to16/N1 ), .Z(
        \pixelfeed/fifo64to16/N84 ) );
  GTECH_NOT \pixelfeed/fifo64to16/I_1  ( .A(\pixelfeed/fifo64to16/produce[0] ), 
        .Z(\pixelfeed/fifo64to16/N0 ) );
  GTECH_AND2 \pixelfeed/fifo64to16/C1682  ( .A(\pixelfeed/fifo64to16/N0 ), .B(
        \pixelfeed/fifo64to16/produce[1] ), .Z(\pixelfeed/fifo64to16/N83 ) );
  GTECH_AND2 \pixelfeed/fifo64to16/C1681  ( .A(
        \pixelfeed/fifo64to16/produce[0] ), .B(
        \pixelfeed/fifo64to16/produce[1] ), .Z(\pixelfeed/fifo64to16/N82 ) );
  SUB_UNS_OP \pixelfeed/fifo64to16/sub_68  ( .A({\pixelfeed/fifo64to16/N38 , 
        \pixelfeed/fifo64to16/N39 , \pixelfeed/fifo64to16/N40 , 
        \pixelfeed/fifo64to16/N41 , \pixelfeed/fifo64to16/N42 }), .B(1'b1), 
        .Z({\pixelfeed/fifo64to16/N52 , \pixelfeed/fifo64to16/N51 , 
        \pixelfeed/fifo64to16/N50 , \pixelfeed/fifo64to16/N49 , 
        \pixelfeed/fifo64to16/N48 }) );
  ADD_UNS_OP \pixelfeed/fifo64to16/add_67  ( .A({
        \pixelfeed/fifo64to16/consume[3] , \pixelfeed/fifo64to16/consume[2] , 
        \pixelfeed/fifo64to16/consume[1] , \pixelfeed/fifo64to16/consume[0] }), 
        .B(1'b1), .Z({\pixelfeed/fifo64to16/N47 , \pixelfeed/fifo64to16/N46 , 
        \pixelfeed/fifo64to16/N45 , \pixelfeed/fifo64to16/N44 }) );
  ADD_UNS_OP \pixelfeed/fifo64to16/add_64  ( .A({
        \pixelfeed/fifo64to16/level[4] , \pixelfeed/fifo64to16/level[3] , 
        \pixelfeed/fifo64to16/level[2] , \pixelfeed/fifo64to16/level[1] , 
        \pixelfeed/fifo64to16/level[0] }), .B({1'b1, 1'b0, 1'b0}), .Z({
        \pixelfeed/fifo64to16/N33 , \pixelfeed/fifo64to16/N32 , 
        \pixelfeed/fifo64to16/N31 , \pixelfeed/fifo64to16/N30 , 
        \pixelfeed/fifo64to16/N29 }) );
  ADD_UNS_OP \pixelfeed/fifo64to16/add_63  ( .A({
        \pixelfeed/fifo64to16/produce[1] , \pixelfeed/fifo64to16/produce[0] }), 
        .B(1'b1), .Z({\pixelfeed/fifo64to16/N28 , \pixelfeed/fifo64to16/N27 })
         );
  GTECH_NOT \pixelfeed/fifo64to16/I_0  ( .A(\pixelfeed/fifo64to16/N80 ), .Z(
        \pixelfeed/fifo64to16/N81 ) );
  GTECH_OR2 \pixelfeed/fifo64to16/C1679  ( .A(\pixelfeed/fifo64to16/level[0] ), 
        .B(\pixelfeed/fifo64to16/N79 ), .Z(\pixelfeed/fifo64to16/N80 ) );
  GTECH_OR2 \pixelfeed/fifo64to16/C1678  ( .A(\pixelfeed/fifo64to16/level[1] ), 
        .B(\pixelfeed/fifo64to16/N78 ), .Z(\pixelfeed/fifo64to16/N79 ) );
  GTECH_OR2 \pixelfeed/fifo64to16/C1677  ( .A(\pixelfeed/fifo64to16/level[2] ), 
        .B(\pixelfeed/fifo64to16/N77 ), .Z(\pixelfeed/fifo64to16/N78 ) );
  GTECH_OR2 \pixelfeed/fifo64to16/C1676  ( .A(\pixelfeed/fifo64to16/level[3] ), 
        .B(\pixelfeed/fifo64to16/level[4] ), .Z(\pixelfeed/fifo64to16/N77 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__0_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__0_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [0]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__1_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__1_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [1]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__2_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__2_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [2]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__3_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__3_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [3]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__4_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__4_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [4]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__5_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__5_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [5]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__6_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__6_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [6]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__7_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__7_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [7]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__8_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__8_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [8]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__9_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__9_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [9]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__10_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__10_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [10]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__11_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__11_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [11]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__12_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__12_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [12]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__13_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__13_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [13]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__14_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__14_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [14]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__15_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__15_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [15]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__16_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__16_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [16]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__17_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__17_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [17]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__18_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__18_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [18]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__19_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__19_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [19]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__20_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__20_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [20]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__21_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__21_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [21]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__22_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__22_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [22]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__23_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__23_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [23]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__24_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__24_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [24]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__25_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__25_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [25]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__26_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__26_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [26]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__27_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__27_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [27]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__28_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__28_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [28]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__29_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__29_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [29]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__30_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__30_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [30]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__31_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__31_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [31]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__32_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__32_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [32]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__33_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__33_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [33]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__34_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__34_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [34]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__35_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__35_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [35]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__36_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__36_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [36]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__37_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__37_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [37]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__38_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__38_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [38]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__39_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__39_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [39]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__40_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__40_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [40]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__41_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__41_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [41]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__42_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__42_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [42]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__43_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__43_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [43]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__44_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__44_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [44]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__45_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__45_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [45]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__46_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__46_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [46]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__47_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__47_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [47]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__48_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__48_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [48]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__49_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__49_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [49]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__50_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__50_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [50]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__51_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__51_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [51]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__52_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__52_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [52]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__53_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__53_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [53]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__54_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__54_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [54]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__55_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__55_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [55]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__56_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__56_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [56]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__57_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__57_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [57]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__58_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__58_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [58]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__59_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__59_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [59]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__60_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__60_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [60]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__61_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__61_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [61]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__62_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__62_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [62]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_3__63_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__63_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [63]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N73 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__0_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__0_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [64]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__1_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__1_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [65]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__2_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__2_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [66]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__3_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__3_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [67]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__4_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__4_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [68]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__5_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__5_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [69]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__6_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__6_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [70]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__7_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__7_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [71]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__8_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__8_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [72]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__9_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__9_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [73]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__10_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__10_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [74]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__11_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__11_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [75]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__12_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__12_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [76]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__13_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__13_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [77]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__14_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__14_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [78]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__15_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__15_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [79]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__16_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__16_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [80]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__17_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__17_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [81]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__18_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__18_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [82]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__19_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__19_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [83]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__20_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__20_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [84]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__21_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__21_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [85]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__22_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__22_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [86]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__23_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__23_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [87]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__24_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__24_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [88]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__25_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__25_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [89]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__26_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__26_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [90]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__27_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__27_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [91]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__28_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__28_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [92]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__29_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__29_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [93]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__30_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__30_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [94]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__31_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__31_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [95]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__32_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__32_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [96]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__33_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__33_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [97]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__34_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__34_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [98]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__35_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__35_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [99]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__36_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__36_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [100]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__37_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__37_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [101]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__38_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__38_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [102]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__39_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__39_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [103]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__40_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__40_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [104]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__41_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__41_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [105]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__42_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__42_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [106]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__43_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__43_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [107]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__44_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__44_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [108]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__45_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__45_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [109]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__46_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__46_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [110]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__47_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__47_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [111]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__48_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__48_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [112]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__49_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__49_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [113]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__50_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__50_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [114]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__51_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__51_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [115]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__52_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__52_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [116]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__53_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__53_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [117]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__54_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__54_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [118]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__55_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__55_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [119]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__56_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__56_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [120]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__57_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__57_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [121]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__58_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__58_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [122]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__59_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__59_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [123]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__60_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__60_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [124]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__61_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__61_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [125]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__62_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__62_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [126]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_2__63_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__63_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [127]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N74 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__0_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__0_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [128]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__1_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__1_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [129]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__2_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__2_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [130]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__3_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__3_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [131]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__4_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__4_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [132]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__5_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__5_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [133]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__6_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__6_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [134]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__7_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__7_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [135]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__8_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__8_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [136]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__9_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__9_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [137]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__10_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__10_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [138]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__11_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__11_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [139]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__12_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__12_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [140]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__13_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__13_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [141]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__14_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__14_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [142]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__15_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__15_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [143]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__16_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__16_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [144]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__17_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__17_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [145]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__18_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__18_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [146]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__19_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__19_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [147]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__20_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__20_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [148]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__21_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__21_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [149]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__22_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__22_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [150]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__23_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__23_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [151]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__24_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__24_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [152]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__25_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__25_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [153]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__26_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__26_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [154]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__27_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__27_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [155]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__28_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__28_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [156]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__29_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__29_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [157]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__30_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__30_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [158]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__31_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__31_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [159]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__32_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__32_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [160]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__33_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__33_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [161]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__34_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__34_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [162]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__35_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__35_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [163]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__36_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__36_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [164]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__37_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__37_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [165]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__38_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__38_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [166]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__39_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__39_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [167]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__40_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__40_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [168]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__41_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__41_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [169]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__42_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__42_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [170]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__43_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__43_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [171]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__44_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__44_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [172]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__45_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__45_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [173]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__46_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__46_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [174]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__47_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__47_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [175]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__48_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__48_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [176]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__49_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__49_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [177]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__50_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__50_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [178]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__51_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__51_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [179]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__52_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__52_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [180]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__53_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__53_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [181]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__54_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__54_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [182]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__55_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__55_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [183]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__56_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__56_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [184]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__57_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__57_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [185]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__58_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__58_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [186]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__59_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__59_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [187]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__60_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__60_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [188]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__61_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__61_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [189]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__62_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__62_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [190]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_1__63_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__63_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [191]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N75 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__0_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__0_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [192]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__1_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__1_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [193]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__2_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__2_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [194]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__3_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__3_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [195]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__4_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__4_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [196]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__5_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__5_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [197]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__6_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__6_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [198]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__7_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__7_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [199]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__8_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__8_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [200]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__9_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__9_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [201]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__10_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__10_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [202]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__11_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__11_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [203]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__12_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__12_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [204]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__13_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__13_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [205]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__14_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__14_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [206]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__15_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__15_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [207]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__16_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__16_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [208]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__17_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__17_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [209]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__18_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__18_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [210]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__19_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__19_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [211]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__20_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__20_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [212]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__21_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__21_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [213]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__22_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__22_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [214]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__23_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__23_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [215]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__24_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__24_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [216]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__25_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__25_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [217]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__26_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__26_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [218]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__27_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__27_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [219]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__28_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__28_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [220]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__29_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__29_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [221]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__30_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__30_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [222]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__31_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__31_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [223]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__32_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__32_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [224]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__33_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__33_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [225]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__34_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__34_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [226]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__35_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__35_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [227]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__36_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__36_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [228]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__37_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__37_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [229]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__38_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__38_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [230]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__39_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__39_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [231]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__40_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__40_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [232]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__41_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__41_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [233]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__42_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__42_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [234]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__43_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__43_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [235]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__44_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__44_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [236]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__45_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__45_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [237]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__46_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__46_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [238]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__47_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__47_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [239]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__48_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__48_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [240]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__49_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__49_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [241]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__50_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__50_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [242]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__51_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__51_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [243]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__52_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__52_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [244]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__53_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__53_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [245]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__54_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__54_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [246]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__55_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__55_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [247]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__56_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__56_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [248]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__57_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__57_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [249]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__58_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__58_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [250]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__59_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__59_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [251]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__60_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__60_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [252]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__61_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__61_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [253]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__62_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__62_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [254]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/storage_reg_0__63_  ( .clear(1'b0), 
        .preset(1'b0), .next_state(\pixelfeed/n_0_net__63_ ), .clocked_on(
        sys_clk), .data_in(1'b0), .enable(1'b0), .Q(
        \pixelfeed/fifo64to16/storage [255]), .QN(), .synch_clear(1'b0), 
        .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        \pixelfeed/fifo64to16/N76 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/consume_reg_0_  ( .clear(1'b0), .preset(
        1'b0), .next_state(\pixelfeed/fifo64to16/N63 ), .clocked_on(sys_clk), 
        .data_in(1'b0), .enable(1'b0), .Q(\pixelfeed/fifo64to16/consume[0] ), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(\pixelfeed/fifo64to16/N62 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/consume_reg_1_  ( .clear(1'b0), .preset(
        1'b0), .next_state(\pixelfeed/fifo64to16/N64 ), .clocked_on(sys_clk), 
        .data_in(1'b0), .enable(1'b0), .Q(\pixelfeed/fifo64to16/consume[1] ), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(\pixelfeed/fifo64to16/N62 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/consume_reg_2_  ( .clear(1'b0), .preset(
        1'b0), .next_state(\pixelfeed/fifo64to16/N65 ), .clocked_on(sys_clk), 
        .data_in(1'b0), .enable(1'b0), .Q(\pixelfeed/fifo64to16/consume[2] ), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(\pixelfeed/fifo64to16/N62 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/consume_reg_3_  ( .clear(1'b0), .preset(
        1'b0), .next_state(\pixelfeed/fifo64to16/N66 ), .clocked_on(sys_clk), 
        .data_in(1'b0), .enable(1'b0), .Q(\pixelfeed/fifo64to16/consume[3] ), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(\pixelfeed/fifo64to16/N62 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/level_reg_0_  ( .clear(1'b0), .preset(
        1'b0), .next_state(\pixelfeed/fifo64to16/N68 ), .clocked_on(sys_clk), 
        .data_in(1'b0), .enable(1'b0), .Q(\pixelfeed/fifo64to16/level[0] ), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(\pixelfeed/fifo64to16/N67 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/level_reg_1_  ( .clear(1'b0), .preset(
        1'b0), .next_state(\pixelfeed/fifo64to16/N69 ), .clocked_on(sys_clk), 
        .data_in(1'b0), .enable(1'b0), .Q(\pixelfeed/fifo64to16/level[1] ), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(\pixelfeed/fifo64to16/N67 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/level_reg_2_  ( .clear(1'b0), .preset(
        1'b0), .next_state(\pixelfeed/fifo64to16/N70 ), .clocked_on(sys_clk), 
        .data_in(1'b0), .enable(1'b0), .Q(\pixelfeed/fifo64to16/level[2] ), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(\pixelfeed/fifo64to16/N67 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/level_reg_3_  ( .clear(1'b0), .preset(
        1'b0), .next_state(\pixelfeed/fifo64to16/N71 ), .clocked_on(sys_clk), 
        .data_in(1'b0), .enable(1'b0), .Q(\pixelfeed/fifo64to16/level[3] ), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(\pixelfeed/fifo64to16/N67 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/level_reg_4_  ( .clear(1'b0), .preset(
        1'b0), .next_state(\pixelfeed/fifo64to16/N72 ), .clocked_on(sys_clk), 
        .data_in(1'b0), .enable(1'b0), .Q(\pixelfeed/fifo64to16/level[4] ), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(\pixelfeed/fifo64to16/N67 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/produce_reg_0_  ( .clear(1'b0), .preset(
        1'b0), .next_state(\pixelfeed/fifo64to16/N60 ), .clocked_on(sys_clk), 
        .data_in(1'b0), .enable(1'b0), .Q(\pixelfeed/fifo64to16/produce[0] ), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(\pixelfeed/fifo64to16/N59 ) );
  \**SEQGEN**  \pixelfeed/fifo64to16/produce_reg_1_  ( .clear(1'b0), .preset(
        1'b0), .next_state(\pixelfeed/fifo64to16/N61 ), .clocked_on(sys_clk), 
        .data_in(1'b0), .enable(1'b0), .Q(\pixelfeed/fifo64to16/produce[1] ), 
        .QN(), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(\pixelfeed/fifo64to16/N59 ) );
  GTECH_AND2 \pixelfeed/fifo64to16/C14  ( .A(\pixelfeed/fifo64to16/consume[1] ), .B(\pixelfeed/fifo64to16/consume[0] ), .Z(\pixelfeed/fifo64to16/N23 ) );
  GTECH_OR2 \pixelfeed/fifo64to16/C12  ( .A(\pixelfeed/fifo64to16/N16 ), .B(
        \pixelfeed/fifo64to16/consume[0] ), .Z(\pixelfeed/fifo64to16/N21 ) );
  GTECH_OR2 \pixelfeed/fifo64to16/C9  ( .A(\pixelfeed/fifo64to16/consume[1] ), 
        .B(\pixelfeed/fifo64to16/N17 ), .Z(\pixelfeed/fifo64to16/N19 ) );
  GTECH_AND2 \pixelfeed/fifo64to16/C7  ( .A(\pixelfeed/fifo64to16/N16 ), .B(
        \pixelfeed/fifo64to16/N17 ), .Z(\pixelfeed/fifo64to16/N18 ) );
endmodule

