
module divider_dshift ( i_clk, i_rst, i_dividend, i_divisor, i_start, o_ready, 
        o_quotient, o_remainder );
  input [31:0] i_dividend;
  input [31:0] i_divisor;
  output [31:0] o_quotient;
  output [31:0] o_remainder;
  input i_clk, i_rst, i_start;
  output o_ready;
  wire   ready, reg_carry, n_1_net__3_, n_1_net__2_, n_1_net__1_, n_1_net__0_,
         state_reg_1_0, N264, N265, N266, N267, N268, N269, N270, N271, N272,
         N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283,
         N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294,
         N295, n701, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n829, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n870, n934, n935, n936, n937, n938, n939, n940, n941, n944,
         n945, n946, n947, n948, n949, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1113, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1296, n1297,
         n1769, n1770, n1771, n1772, n1773, n1864, n1988, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, \shifter_0/n49 , \shifter_0/n48 ,
         \shifter_0/n47 , \shifter_0/n46 , \shifter_0/n45 , \shifter_0/n44 ,
         \shifter_0/n43 , \shifter_0/n42 , \shifter_0/n41 , \shifter_0/n40 ,
         \shifter_0/n39 , \shifter_0/n38 , \shifter_0/n37 , \shifter_0/n36 ,
         \shifter_0/n35 , \shifter_0/n34 , \shifter_0/n33 , \shifter_0/n32 ,
         \shifter_0/n31 , \shifter_0/n30 , \shifter_0/o_shifted[4] ,
         \shifter_0/n20 , \shifter_0/n4 , \shifter_0/n3 , \shifter_0/n2 ,
         \shifter_0/n1 , \shifter_0/n25 , \shifter_0/n24 , \shifter_0/n21 ,
         \shifter_0/shift_1b_0/n33 , \shifter_0/shift_3b_0/n38 ,
         \shifter_0/shift_3b_0/n37 , \shifter_0/shift_3b_0/n36 ,
         \shifter_0/shift_3b_0/n35 , \shifter_0/shift_3b_0/n13 ,
         \shifter_0/shift_3b_0/n5 , \shifter_0/shift_3b_0/n4 ,
         \shifter_0/shift_3b_0/n3 , \shifter_0/shift_3b_0/n2 ,
         \shifter_0/shift_3b_0/n34 , \shifter_0/shift_3b_0/n33 ,
         \shifter_0/shift_3b_0/n32 , \shifter_0/shift_3b_0/n31 ,
         \shifter_0/shift_3b_0/n30 , \shifter_0/shift_3b_0/n29 ,
         \shifter_0/shift_3b_0/n28 , \shifter_0/shift_3b_0/n27 ,
         \shifter_0/shift_3b_0/n26 , \shifter_0/shift_3b_0/n25 ,
         \shifter_0/shift_3b_0/n24 , \shifter_0/shift_3b_0/n23 ,
         \shifter_0/shift_3b_0/n22 , \shifter_0/shift_3b_0/n21 ,
         \shifter_0/shift_3b_0/n20 , \shifter_0/shift_3b_0/n19 ,
         \shifter_0/shift_3b_0/n18 , \shifter_0/shift_3b_0/n14 ,
         \shifter_0/shift_3b_0/n12 , \shifter_0/shift_3b_0/n11 ,
         \shifter_0/shift_3b_0/n10 , \shifter_0/shift_3b_0/n9 ,
         \shifter_0/shift_3b_0/n8 , \shifter_0/shift_3b_0/n7 ,
         \shifter_0/shift_3b_0/n6 , \shifter_0/shift_3b_0/shift1 ,
         \shifter_0/shift_3b_0/shift_1b_0/n33 , \shifter_0/shift_3b_1/n38 ,
         \shifter_0/shift_3b_1/n37 , \shifter_0/shift_3b_1/n36 ,
         \shifter_0/shift_3b_1/n35 , \shifter_0/shift_3b_1/n14 ,
         \shifter_0/shift_3b_1/n4 , \shifter_0/shift_3b_1/n3 ,
         \shifter_0/shift_3b_1/n2 , \shifter_0/shift_3b_1/n34 ,
         \shifter_0/shift_3b_1/n33 , \shifter_0/shift_3b_1/n32 ,
         \shifter_0/shift_3b_1/n31 , \shifter_0/shift_3b_1/n30 ,
         \shifter_0/shift_3b_1/n29 , \shifter_0/shift_3b_1/n28 ,
         \shifter_0/shift_3b_1/n27 , \shifter_0/shift_3b_1/n26 ,
         \shifter_0/shift_3b_1/n25 , \shifter_0/shift_3b_1/n24 ,
         \shifter_0/shift_3b_1/n23 , \shifter_0/shift_3b_1/n22 ,
         \shifter_0/shift_3b_1/n21 , \shifter_0/shift_3b_1/n20 ,
         \shifter_0/shift_3b_1/n19 , \shifter_0/shift_3b_1/n16 ,
         \shifter_0/shift_3b_1/n13 , \shifter_0/shift_3b_1/n12 ,
         \shifter_0/shift_3b_1/n11 , \shifter_0/shift_3b_1/n10 ,
         \shifter_0/shift_3b_1/n9 , \shifter_0/shift_3b_1/n8 ,
         \shifter_0/shift_3b_1/n7 , \shifter_0/shift_3b_1/n6 ,
         \shifter_0/shift_3b_1/n5 , \shifter_0/shift_3b_1/shift1 ,
         \shifter_0/shift_3b_1/shift_1b_0/n33 , \shifter_0/shift_7b_0/n48 ,
         \shifter_0/shift_7b_0/n47 , \shifter_0/shift_7b_0/n46 ,
         \shifter_0/shift_7b_0/n45 , \shifter_0/shift_7b_0/n44 ,
         \shifter_0/shift_7b_0/n43 , \shifter_0/shift_7b_0/n42 ,
         \shifter_0/shift_7b_0/n41 , \shifter_0/shift_7b_0/n40 ,
         \shifter_0/shift_7b_0/n39 , \shifter_0/shift_7b_0/n21 ,
         \shifter_0/shift_7b_0/n10 , \shifter_0/shift_7b_0/n9 ,
         \shifter_0/shift_7b_0/n8 , \shifter_0/shift_7b_0/n7 ,
         \shifter_0/shift_7b_0/n6 , \shifter_0/shift_7b_0/n5 ,
         \shifter_0/shift_7b_0/n4 , \shifter_0/shift_7b_0/n38 ,
         \shifter_0/shift_7b_0/n37 , \shifter_0/shift_7b_0/n36 ,
         \shifter_0/shift_7b_0/n35 , \shifter_0/shift_7b_0/n34 ,
         \shifter_0/shift_7b_0/n33 , \shifter_0/shift_7b_0/n32 ,
         \shifter_0/shift_7b_0/n31 , \shifter_0/shift_7b_0/n30 ,
         \shifter_0/shift_7b_0/n29 , \shifter_0/shift_7b_0/n20 ,
         \shifter_0/shift_7b_0/n19 , \shifter_0/shift_7b_0/n18 ,
         \shifter_0/shift_7b_0/n17 , \shifter_0/shift_7b_0/n16 ,
         \shifter_0/shift_7b_0/n15 , \shifter_0/shift_7b_0/n14 ,
         \shifter_0/shift_7b_0/n13 , \shifter_0/shift_7b_0/n12 ,
         \shifter_0/shift_7b_0/n11 , \shifter_0/shift_7b_0/shift_3b_0/n38 ,
         \shifter_0/shift_7b_0/shift_3b_0/n37 ,
         \shifter_0/shift_7b_0/shift_3b_0/n36 ,
         \shifter_0/shift_7b_0/shift_3b_0/n35 ,
         \shifter_0/shift_7b_0/shift_3b_0/n18 ,
         \shifter_0/shift_7b_0/shift_3b_0/n4 ,
         \shifter_0/shift_7b_0/shift_3b_0/n3 ,
         \shifter_0/shift_7b_0/shift_3b_0/n2 ,
         \shifter_0/shift_7b_0/shift_3b_0/n34 ,
         \shifter_0/shift_7b_0/shift_3b_0/n33 ,
         \shifter_0/shift_7b_0/shift_3b_0/n32 ,
         \shifter_0/shift_7b_0/shift_3b_0/n31 ,
         \shifter_0/shift_7b_0/shift_3b_0/n30 ,
         \shifter_0/shift_7b_0/shift_3b_0/n29 ,
         \shifter_0/shift_7b_0/shift_3b_0/n28 ,
         \shifter_0/shift_7b_0/shift_3b_0/n27 ,
         \shifter_0/shift_7b_0/shift_3b_0/n26 ,
         \shifter_0/shift_7b_0/shift_3b_0/n25 ,
         \shifter_0/shift_7b_0/shift_3b_0/n24 ,
         \shifter_0/shift_7b_0/shift_3b_0/n23 ,
         \shifter_0/shift_7b_0/shift_3b_0/n20 ,
         \shifter_0/shift_7b_0/shift_3b_0/n17 ,
         \shifter_0/shift_7b_0/shift_3b_0/n16 ,
         \shifter_0/shift_7b_0/shift_3b_0/n15 ,
         \shifter_0/shift_7b_0/shift_3b_0/n14 ,
         \shifter_0/shift_7b_0/shift_3b_0/n13 ,
         \shifter_0/shift_7b_0/shift_3b_0/n12 ,
         \shifter_0/shift_7b_0/shift_3b_0/n11 ,
         \shifter_0/shift_7b_0/shift_3b_0/n10 ,
         \shifter_0/shift_7b_0/shift_3b_0/n9 ,
         \shifter_0/shift_7b_0/shift_3b_0/n8 ,
         \shifter_0/shift_7b_0/shift_3b_0/n7 ,
         \shifter_0/shift_7b_0/shift_3b_0/n6 ,
         \shifter_0/shift_7b_0/shift_3b_0/n5 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift1 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n33 , \adder_0/G6_1 ,
         \adder_0/G6_3 , \adder_0/G6_5 , \adder_0/G6_7 , \adder_0/G6_9 ,
         \adder_0/G6_11 , \adder_0/G6_13 , \adder_0/G6_15 , \adder_0/G6_17 ,
         \adder_0/G6_19 , \adder_0/G6_21 , \adder_0/G6_23 , \adder_0/G6_25 ,
         \adder_0/G6_27 , \adder_0/G6_29_ , \adder_0/G5[8] , \adder_0/G5[9] ,
         \adder_0/G5[10] , \adder_0/G5[11] , \adder_0/G5[12] ,
         \adder_0/G5[13] , \adder_0/G5[14] , \adder_0/G5[15] , \adder_0/G4[4] ,
         \adder_0/G4[5] , \adder_0/G4[6] , \adder_0/G4[7] , \adder_0/G4[8] ,
         \adder_0/G4[9] , \adder_0/G4[10] , \adder_0/G4[11] , \adder_0/G4[12] ,
         \adder_0/G4[13] , \adder_0/G4[14] , \adder_0/G4[15] , \adder_0/P3[4] ,
         \adder_0/P3[5] , \adder_0/P3[6] , \adder_0/P3[7] , \adder_0/P3[8] ,
         \adder_0/P3[9] , \adder_0/P3[10] , \adder_0/P3[11] , \adder_0/P3[12] ,
         \adder_0/P3[13] , \adder_0/P3[14] , \adder_0/P3[15] , \adder_0/G3[2] ,
         \adder_0/G3[3] , \adder_0/G3[4] , \adder_0/G3[5] , \adder_0/G3[6] ,
         \adder_0/G3[7] , \adder_0/G3[8] , \adder_0/G3[9] , \adder_0/G3[10] ,
         \adder_0/G3[11] , \adder_0/G3[12] , \adder_0/G3[13] ,
         \adder_0/G3[14] , \adder_0/G3[15] , \adder_0/P2[2] , \adder_0/P2[3] ,
         \adder_0/P2[4] , \adder_0/P2[5] , \adder_0/P2[6] , \adder_0/P2[7] ,
         \adder_0/P2[8] , \adder_0/P2[9] , \adder_0/P2[10] , \adder_0/P2[11] ,
         \adder_0/P2[12] , \adder_0/P2[13] , \adder_0/P2[14] ,
         \adder_0/P2[15] , \adder_0/G2[1] , \adder_0/G2[2] , \adder_0/G2[3] ,
         \adder_0/G2[4] , \adder_0/G2[5] , \adder_0/G2[6] , \adder_0/G2[7] ,
         \adder_0/G2[8] , \adder_0/G2[9] , \adder_0/G2[10] , \adder_0/G2[11] ,
         \adder_0/G2[12] , \adder_0/G2[13] , \adder_0/G2[14] ,
         \adder_0/G2[15] , \adder_0/P1[1] , \adder_0/P1[2] , \adder_0/P1[3] ,
         \adder_0/P1[4] , \adder_0/P1[5] , \adder_0/P1[6] , \adder_0/P1[7] ,
         \adder_0/P1[8] , \adder_0/P1[9] , \adder_0/P1[10] , \adder_0/P1[11] ,
         \adder_0/P1[12] , \adder_0/P1[13] , \adder_0/P1[14] ,
         \adder_0/P1[15] , \adder_0/G1[0] , \adder_0/G1[1] , \adder_0/G1[2] ,
         \adder_0/G1[3] , \adder_0/G1[4] , \adder_0/G1[5] , \adder_0/G1[6] ,
         \adder_0/G1[7] , \adder_0/G1[8] , \adder_0/G1[9] , \adder_0/G1[10] ,
         \adder_0/G1[11] , \adder_0/G1[12] , \adder_0/G1[13] ,
         \adder_0/G1[14] , \adder_0/G1[15] , \adder_0/G0[0] , \adder_0/G0[1] ,
         \adder_0/G0[2] , \adder_0/G0[3] , \adder_0/G0[4] , \adder_0/G0[5] ,
         \adder_0/G0[6] , \adder_0/G0[7] , \adder_0/G0[8] , \adder_0/G0[9] ,
         \adder_0/G0[10] , \adder_0/G0[11] , \adder_0/G0[12] ,
         \adder_0/G0[13] , \adder_0/G0[14] , \adder_0/G0[15] ,
         \adder_0/G0[16] , \adder_0/G0[17] , \adder_0/G0[18] ,
         \adder_0/G0[19] , \adder_0/G0[20] , \adder_0/G0[21] ,
         \adder_0/G0[22] , \adder_0/G0[23] , \adder_0/G0[24] ,
         \adder_0/G0[25] , \adder_0/G0[26] , \adder_0/G0[27] ,
         \adder_0/G0[28] , \adder_0/G0[29] , \adder_0/G0[30] ,
         \adder_0/G0[31] , \adder_0/P0[0] , \adder_0/P0[1] , \adder_0/P0[2] ,
         \adder_0/P0[3] , \adder_0/P0[4] , \adder_0/P0[5] , \adder_0/P0[6] ,
         \adder_0/P0[7] , \adder_0/P0[8] , \adder_0/P0[9] , \adder_0/P0[10] ,
         \adder_0/P0[11] , \adder_0/P0[12] , \adder_0/P0[13] ,
         \adder_0/P0[14] , \adder_0/P0[15] , \adder_0/P0[16] ,
         \adder_0/P0[17] , \adder_0/P0[18] , \adder_0/P0[19] ,
         \adder_0/P0[20] , \adder_0/P0[21] , \adder_0/P0[22] ,
         \adder_0/P0[23] , \adder_0/P0[24] , \adder_0/P0[25] ,
         \adder_0/P0[26] , \adder_0/P0[27] , \adder_0/P0[28] ,
         \adder_0/P0[29] , \adder_0/P0[30] , \adder_0/P0[31] , \adder_0/o_c ,
         \adder_0/operator_C_stage_1_0/n3 , \adder_0/operator_B_stage_1_1/n3 ,
         \adder_0/operator_B_stage_1_2/n3 , \adder_0/operator_B_stage_1_3/n3 ,
         \adder_0/operator_B_stage_1_4/n3 , \adder_0/operator_B_stage_1_5/n3 ,
         \adder_0/operator_B_stage_1_6/n3 , \adder_0/operator_B_stage_1_7/n3 ,
         \adder_0/operator_B_stage_1_8/n3 , \adder_0/operator_B_stage_1_9/n3 ,
         \adder_0/operator_B_stage_1_10/n3 ,
         \adder_0/operator_B_stage_1_11/n3 ,
         \adder_0/operator_B_stage_1_12/n3 ,
         \adder_0/operator_B_stage_1_13/n3 ,
         \adder_0/operator_B_stage_1_14/n3 ,
         \adder_0/operator_B_stage_1_15/n3 , \adder_0/operator_C_stage_2_1/n3 ,
         \adder_0/operator_B_stage_2_2/n3 , \adder_0/operator_B_stage_2_3/n3 ,
         \adder_0/operator_B_stage_2_4/n3 , \adder_0/operator_B_stage_2_5/n3 ,
         \adder_0/operator_B_stage_2_6/n3 , \adder_0/operator_B_stage_2_7/n3 ,
         \adder_0/operator_B_stage_2_8/n3 , \adder_0/operator_B_stage_2_9/n3 ,
         \adder_0/operator_B_stage_2_10/n3 ,
         \adder_0/operator_B_stage_2_11/n3 ,
         \adder_0/operator_B_stage_2_12/n3 ,
         \adder_0/operator_B_stage_2_13/n3 ,
         \adder_0/operator_B_stage_2_14/n3 ,
         \adder_0/operator_B_stage_2_15/n3 , \adder_0/operator_C_stage_3_2/n3 ,
         \adder_0/operator_C_stage_3_3/n3 , \adder_0/operator_B_stage_3_4/n3 ,
         \adder_0/operator_B_stage_3_5/n3 , \adder_0/operator_B_stage_3_6/n3 ,
         \adder_0/operator_B_stage_3_7/n3 , \adder_0/operator_B_stage_3_8/n3 ,
         \adder_0/operator_B_stage_3_9/n3 , \adder_0/operator_B_stage_3_10/n3 ,
         \adder_0/operator_B_stage_3_11/n3 ,
         \adder_0/operator_B_stage_3_12/n3 ,
         \adder_0/operator_B_stage_3_13/n3 ,
         \adder_0/operator_B_stage_3_14/n3 ,
         \adder_0/operator_B_stage_3_15/n3 , \adder_0/operator_C_stage_4_4/n3 ,
         \adder_0/operator_C_stage_4_5/n3 , \adder_0/operator_C_stage_4_6/n3 ,
         \adder_0/operator_C_stage_4_7/n3 , \adder_0/operator_B_stage_4_8/n3 ,
         \adder_0/operator_B_stage_4_9/n3 , \adder_0/operator_B_stage_4_10/n3 ,
         \adder_0/operator_B_stage_4_11/n3 ,
         \adder_0/operator_B_stage_4_12/n3 ,
         \adder_0/operator_B_stage_4_13/n3 ,
         \adder_0/operator_B_stage_4_14/n3 ,
         \adder_0/operator_B_stage_4_15/n3 , \adder_0/operator_C_stage_5_8/n3 ,
         \adder_0/operator_C_stage_5_9/n3 , \adder_0/operator_C_stage_5_10/n3 ,
         \adder_0/operator_C_stage_5_11/n3 ,
         \adder_0/operator_C_stage_5_12/n3 ,
         \adder_0/operator_C_stage_5_13/n3 ,
         \adder_0/operator_C_stage_5_14/n3 ,
         \adder_0/operator_C_stage_5_15/n3 , \adder_0/operator_C_stage_6_0/n3 ,
         \adder_0/operator_C_stage_6_1/n3 , \adder_0/operator_C_stage_6_2/n3 ,
         \adder_0/operator_C_stage_6_3/n3 , \adder_0/operator_C_stage_6_4/n3 ,
         \adder_0/operator_C_stage_6_5/n3 , \adder_0/operator_C_stage_6_6/n3 ,
         \adder_0/operator_C_stage_6_7/n3 , \adder_0/operator_C_stage_6_8/n3 ,
         \adder_0/operator_C_stage_6_9/n3 , \adder_0/operator_C_stage_6_10/n3 ,
         \adder_0/operator_C_stage_6_11/n3 ,
         \adder_0/operator_C_stage_6_12/n3 ,
         \adder_0/operator_C_stage_6_13/n3 ,
         \adder_0/operator_C_stage_6_14/n3 ,
         \adder_0/operator_C_stage_6_15/n3 , \adder_1/G6_1 , \adder_1/G6_3 ,
         \adder_1/G6_5 , \adder_1/G6_7 , \adder_1/G6_9 , \adder_1/G6_11 ,
         \adder_1/G6_13 , \adder_1/G6_15 , \adder_1/G6_17 , \adder_1/G6_19 ,
         \adder_1/G6_21 , \adder_1/G6_23 , \adder_1/G6_25 , \adder_1/G6_27 ,
         \adder_1/G6_29_ , \adder_1/G5[8] , \adder_1/G5[9] , \adder_1/G5[10] ,
         \adder_1/G5[11] , \adder_1/G5[12] , \adder_1/G5[13] ,
         \adder_1/G5[14] , \adder_1/G5[15] , \adder_1/G4[4] , \adder_1/G4[5] ,
         \adder_1/G4[6] , \adder_1/G4[7] , \adder_1/G4[8] , \adder_1/G4[9] ,
         \adder_1/G4[10] , \adder_1/G4[11] , \adder_1/G4[12] ,
         \adder_1/G4[13] , \adder_1/G4[14] , \adder_1/G4[15] , \adder_1/P3[4] ,
         \adder_1/P3[5] , \adder_1/P3[6] , \adder_1/P3[7] , \adder_1/P3[8] ,
         \adder_1/P3[9] , \adder_1/P3[10] , \adder_1/P3[11] , \adder_1/P3[12] ,
         \adder_1/P3[13] , \adder_1/P3[14] , \adder_1/P3[15] , \adder_1/G3[2] ,
         \adder_1/G3[3] , \adder_1/G3[4] , \adder_1/G3[5] , \adder_1/G3[6] ,
         \adder_1/G3[7] , \adder_1/G3[8] , \adder_1/G3[9] , \adder_1/G3[10] ,
         \adder_1/G3[11] , \adder_1/G3[12] , \adder_1/G3[13] ,
         \adder_1/G3[14] , \adder_1/G3[15] , \adder_1/P2[2] , \adder_1/P2[3] ,
         \adder_1/P2[4] , \adder_1/P2[5] , \adder_1/P2[6] , \adder_1/P2[7] ,
         \adder_1/P2[8] , \adder_1/P2[9] , \adder_1/P2[10] , \adder_1/P2[11] ,
         \adder_1/P2[12] , \adder_1/P2[13] , \adder_1/P2[14] ,
         \adder_1/P2[15] , \adder_1/G2[1] , \adder_1/G2[2] , \adder_1/G2[3] ,
         \adder_1/G2[4] , \adder_1/G2[5] , \adder_1/G2[6] , \adder_1/G2[7] ,
         \adder_1/G2[8] , \adder_1/G2[9] , \adder_1/G2[10] , \adder_1/G2[11] ,
         \adder_1/G2[12] , \adder_1/G2[13] , \adder_1/G2[14] ,
         \adder_1/G2[15] , \adder_1/P1[1] , \adder_1/P1[2] , \adder_1/P1[3] ,
         \adder_1/P1[4] , \adder_1/P1[5] , \adder_1/P1[6] , \adder_1/P1[7] ,
         \adder_1/P1[8] , \adder_1/P1[9] , \adder_1/P1[10] , \adder_1/P1[11] ,
         \adder_1/P1[12] , \adder_1/P1[13] , \adder_1/P1[14] ,
         \adder_1/P1[15] , \adder_1/G1[0] , \adder_1/G1[1] , \adder_1/G1[2] ,
         \adder_1/G1[3] , \adder_1/G1[4] , \adder_1/G1[5] , \adder_1/G1[6] ,
         \adder_1/G1[7] , \adder_1/G1[8] , \adder_1/G1[9] , \adder_1/G1[10] ,
         \adder_1/G1[11] , \adder_1/G1[12] , \adder_1/G1[13] ,
         \adder_1/G1[14] , \adder_1/G1[15] , \adder_1/G0[0] , \adder_1/G0[1] ,
         \adder_1/G0[2] , \adder_1/G0[3] , \adder_1/G0[4] , \adder_1/G0[5] ,
         \adder_1/G0[6] , \adder_1/G0[7] , \adder_1/G0[8] , \adder_1/G0[9] ,
         \adder_1/G0[10] , \adder_1/G0[11] , \adder_1/G0[12] ,
         \adder_1/G0[13] , \adder_1/G0[14] , \adder_1/G0[15] ,
         \adder_1/G0[16] , \adder_1/G0[17] , \adder_1/G0[18] ,
         \adder_1/G0[19] , \adder_1/G0[20] , \adder_1/G0[21] ,
         \adder_1/G0[22] , \adder_1/G0[23] , \adder_1/G0[24] ,
         \adder_1/G0[25] , \adder_1/G0[26] , \adder_1/G0[27] ,
         \adder_1/G0[28] , \adder_1/G0[29] , \adder_1/G0[30] ,
         \adder_1/G0[31] , \adder_1/P0[0] , \adder_1/P0[1] , \adder_1/P0[2] ,
         \adder_1/P0[3] , \adder_1/P0[4] , \adder_1/P0[5] , \adder_1/P0[6] ,
         \adder_1/P0[7] , \adder_1/P0[8] , \adder_1/P0[9] , \adder_1/P0[10] ,
         \adder_1/P0[11] , \adder_1/P0[12] , \adder_1/P0[13] ,
         \adder_1/P0[14] , \adder_1/P0[15] , \adder_1/P0[16] ,
         \adder_1/P0[17] , \adder_1/P0[18] , \adder_1/P0[19] ,
         \adder_1/P0[20] , \adder_1/P0[21] , \adder_1/P0[22] ,
         \adder_1/P0[23] , \adder_1/P0[24] , \adder_1/P0[25] ,
         \adder_1/P0[26] , \adder_1/P0[27] , \adder_1/P0[28] ,
         \adder_1/P0[29] , \adder_1/P0[30] , \adder_1/P0[31] , \adder_1/o_c ,
         \adder_1/operator_C_stage_1_0/n3 , \adder_1/operator_B_stage_1_1/n3 ,
         \adder_1/operator_B_stage_1_2/n3 , \adder_1/operator_B_stage_1_3/n3 ,
         \adder_1/operator_B_stage_1_4/n3 , \adder_1/operator_B_stage_1_5/n3 ,
         \adder_1/operator_B_stage_1_6/n3 , \adder_1/operator_B_stage_1_7/n3 ,
         \adder_1/operator_B_stage_1_8/n3 , \adder_1/operator_B_stage_1_9/n3 ,
         \adder_1/operator_B_stage_1_10/n3 ,
         \adder_1/operator_B_stage_1_11/n3 ,
         \adder_1/operator_B_stage_1_12/n3 ,
         \adder_1/operator_B_stage_1_13/n3 ,
         \adder_1/operator_B_stage_1_14/n3 ,
         \adder_1/operator_B_stage_1_15/n3 , \adder_1/operator_C_stage_2_1/n3 ,
         \adder_1/operator_B_stage_2_2/n3 , \adder_1/operator_B_stage_2_3/n3 ,
         \adder_1/operator_B_stage_2_4/n3 , \adder_1/operator_B_stage_2_5/n3 ,
         \adder_1/operator_B_stage_2_6/n3 , \adder_1/operator_B_stage_2_7/n3 ,
         \adder_1/operator_B_stage_2_8/n3 , \adder_1/operator_B_stage_2_9/n3 ,
         \adder_1/operator_B_stage_2_10/n3 ,
         \adder_1/operator_B_stage_2_11/n3 ,
         \adder_1/operator_B_stage_2_12/n3 ,
         \adder_1/operator_B_stage_2_13/n3 ,
         \adder_1/operator_B_stage_2_14/n3 ,
         \adder_1/operator_B_stage_2_15/n3 , \adder_1/operator_C_stage_3_2/n3 ,
         \adder_1/operator_C_stage_3_3/n3 , \adder_1/operator_B_stage_3_4/n3 ,
         \adder_1/operator_B_stage_3_5/n3 , \adder_1/operator_B_stage_3_6/n3 ,
         \adder_1/operator_B_stage_3_7/n3 , \adder_1/operator_B_stage_3_8/n3 ,
         \adder_1/operator_B_stage_3_9/n3 , \adder_1/operator_B_stage_3_10/n3 ,
         \adder_1/operator_B_stage_3_11/n3 ,
         \adder_1/operator_B_stage_3_12/n3 ,
         \adder_1/operator_B_stage_3_13/n3 ,
         \adder_1/operator_B_stage_3_14/n3 ,
         \adder_1/operator_B_stage_3_15/n3 , \adder_1/operator_C_stage_4_4/n3 ,
         \adder_1/operator_C_stage_4_5/n3 , \adder_1/operator_C_stage_4_6/n3 ,
         \adder_1/operator_C_stage_4_7/n3 , \adder_1/operator_B_stage_4_8/n3 ,
         \adder_1/operator_B_stage_4_9/n3 , \adder_1/operator_B_stage_4_10/n3 ,
         \adder_1/operator_B_stage_4_11/n3 ,
         \adder_1/operator_B_stage_4_12/n3 ,
         \adder_1/operator_B_stage_4_13/n3 ,
         \adder_1/operator_B_stage_4_14/n3 ,
         \adder_1/operator_B_stage_4_15/n3 , \adder_1/operator_C_stage_5_8/n3 ,
         \adder_1/operator_C_stage_5_9/n3 , \adder_1/operator_C_stage_5_10/n3 ,
         \adder_1/operator_C_stage_5_11/n3 ,
         \adder_1/operator_C_stage_5_12/n3 ,
         \adder_1/operator_C_stage_5_13/n3 ,
         \adder_1/operator_C_stage_5_14/n3 ,
         \adder_1/operator_C_stage_5_15/n3 , \adder_1/operator_C_stage_6_0/n3 ,
         \adder_1/operator_C_stage_6_1/n3 , \adder_1/operator_C_stage_6_2/n3 ,
         \adder_1/operator_C_stage_6_3/n3 , \adder_1/operator_C_stage_6_4/n3 ,
         \adder_1/operator_C_stage_6_5/n3 , \adder_1/operator_C_stage_6_6/n3 ,
         \adder_1/operator_C_stage_6_7/n3 , \adder_1/operator_C_stage_6_8/n3 ,
         \adder_1/operator_C_stage_6_9/n3 , \adder_1/operator_C_stage_6_10/n3 ,
         \adder_1/operator_C_stage_6_11/n3 ,
         \adder_1/operator_C_stage_6_12/n3 ,
         \adder_1/operator_C_stage_6_13/n3 ,
         \adder_1/operator_C_stage_6_14/n3 ,
         \adder_1/operator_C_stage_6_15/n3 , \sra_198/n285 , \sra_198/n284 ,
         \sra_198/n283 , \sra_198/n282 , \sra_198/n281 , \sra_198/n280 ,
         \sra_198/n279 , \sra_198/n278 , \sra_198/n277 , \sra_198/n276 ,
         \sra_198/n275 , \sra_198/n274 , \sra_198/n273 , \sra_198/n272 ,
         \sra_198/n271 , \sra_198/n270 , \sra_198/n269 , \sra_198/n268 ,
         \sra_198/n267 , \sra_198/n266 , \sra_198/n265 , \sra_198/n264 ,
         \sra_198/n263 , \sra_198/n262 , \sra_198/n261 , \sra_198/n260 ,
         \sra_198/n259 , \sra_198/n258 , \sra_198/n257 , \sra_198/n256 ,
         \sra_198/n255 , \sra_198/n254 , \sra_198/n253 , \sra_198/n252 ,
         \sra_198/n251 , \sra_198/n250 , \sra_198/n249 , \sra_198/n248 ,
         \sra_198/n247 , \sra_198/n246 , \sra_198/n245 , \sra_198/n244 ,
         \sra_198/n243 , \sra_198/n242 , \sra_198/n241 , \sra_198/n240 ,
         \sra_198/n239 , \sra_198/n238 , \sra_198/n237 , \sra_198/n236 ,
         \sra_198/n235 , \sra_198/n234 , \sra_198/n233 , \sra_198/n232 ,
         \sra_198/n231 , \sra_198/n230 , \sra_198/n229 , \sra_198/n228 ,
         \sra_198/n227 , \sra_198/n226 , \sra_198/n225 , \sra_198/n224 ,
         \sra_198/n223 , \sra_198/n222 , \sra_198/n221 , \sra_198/n220 ,
         \sra_198/n219 , \sra_198/n218 , \sra_198/n217 , \sra_198/n216 ,
         \sra_198/n215 , \sra_198/n214 , \sra_198/n212 , \sra_198/n211 ,
         \sra_198/n210 , \sra_198/n209 , \sra_198/n208 , \sra_198/n207 ,
         \sra_198/n206 , \sra_198/n205 , \sra_198/n204 , \sra_198/n203 ,
         \sra_198/n202 , \sra_198/n201 , \sra_198/n200 , \sra_198/n199 ,
         \sra_198/n198 , \sra_198/n197 , \sra_198/n196 , \sra_198/n195 ,
         \sra_198/n194 , \sra_198/n193 , \sra_198/n192 , \sra_198/n191 ,
         \sra_198/n190 , \sra_198/n189 , \sra_198/n188 , \sra_198/n187 ,
         \sra_198/n186 , \sra_198/n185 , \sra_198/n184 , \sra_198/n183 ,
         \sra_198/n182 , \sra_198/n181 , \sra_198/n180 , \sra_198/n179 ,
         \sra_198/n178 , \sra_198/n177 , \sra_198/n176 , \sra_198/n175 ,
         \sra_198/n174 , \sra_198/n173 , \sra_198/n172 , \sra_198/n171 ,
         \sra_198/n170 , \sra_198/n169 , \sra_198/n168 , \sra_198/n167 ,
         \sra_198/n166 , \sra_198/n165 , \sra_198/n164 , \sra_198/n163 ,
         \sra_198/n162 , \sra_198/n161 , \sra_198/n160 , \sra_198/n159 ,
         \sra_198/n158 , \sra_198/n157 , \sra_198/n156 , \sra_198/n155 ,
         \sra_198/n154 , \sra_198/n153 , \sra_198/n152 , \sra_198/n151 ,
         \sra_198/n150 , \sra_198/n149 , \sra_198/n148 , \sra_198/n147 ,
         \sra_198/n146 , \sra_198/n145 , \sra_198/n144 , \sra_198/n143 ,
         \sra_198/n142 , \sra_198/n141 , \sra_198/n140 , \sra_198/n139 ,
         \sra_198/n138 , \sra_198/n137 , \sra_198/n136 , \sra_198/n135 ,
         \sra_198/n134 , \sra_198/n133 , \sra_198/n132 , \sra_198/n131 ,
         \sra_198/n130 , \sra_198/n129 , \sra_198/n128 , \sra_198/n127 ,
         \sra_198/n126 , \sra_198/n125 , \sra_198/n124 , \sra_198/n123 ,
         \sra_198/n122 , \sra_198/n121 , \sra_198/n120 , \sra_198/n119 ,
         \sra_198/n118 , \sra_198/n117 , \sra_198/n116 , \sra_198/n115 ,
         \sra_198/n114 , \sra_198/n113 , \sra_198/n112 , \sra_198/n111 ,
         \sra_198/n110 , \sra_198/n109 , \sra_198/n108 , \sra_198/n107 ,
         \sra_198/n106 , \sra_198/n105 , \sra_198/n104 , \sra_198/n103 ,
         \sra_198/n102 , \sra_198/n101 , \sra_198/n100 , \sra_198/n99 ,
         \sra_198/n98 , \sra_198/n97 , \sra_198/n96 , \sra_198/n95 ,
         \sra_198/n94 , \sra_198/n93 , \sra_198/n92 , \sra_198/n91 ,
         \sra_198/n90 , \sra_198/n89 , \sra_198/n88 , \sra_198/n87 ,
         \sra_198/n86 , \sra_198/n85 , \sra_198/n84 , \sra_198/n83 ,
         \sra_198/n82 , \sra_198/n81 , \sra_198/n80 , \sra_198/n79 ,
         \sra_198/n78 , \sra_198/n77 , \sra_198/n76 , \sra_198/n75 ,
         \sra_198/n74 ;
  wire   [30:0] nq;
  wire   [30:0] nqp1;
  wire   [30:0] q;
  wire   [30:0] qp1;
  wire   [31:0] sdata;
  wire   [31:0] sdata_o;
  wire   [3:0] shifted_o;
  wire   [5:0] state;
  wire   [5:0] ct_1;
  wire   [31:0] PR_1;
  wire   [31:0] reg_a;
  wire   [31:0] reg_b;
  wire   [31:0] sum;
  wire   [5:0] sum_ct;
  wire   [5:0] ct;
  wire   [31:0] \shifter_0/data_3 ;
  wire   [31:0] \shifter_0/data_2 ;
  wire   [31:0] \shifter_0/data_1 ;
  wire   [1:0] \shifter_0/shift_3b_0/data1 ;
  wire   [1:0] \shifter_0/shift_3b_1/data1 ;
  wire   [2:0] \shifter_0/shift_7b_0/shift1 ;
  wire   [3:0] \shifter_0/shift_7b_0/data1 ;
  wire   [1:0] \shifter_0/shift_7b_0/shift_3b_0/data1 ;
  wire   [15:8] \adder_0/P4 ;
  wire   [15:8] \adder_1/P4 ;
  wire   [30:2] \add_35/carry ;
  wire   [30:2] \add_34/carry ;

  DFFR_X1 PR_reg_0_ ( .D(n3355), .CK(i_clk), .RN(i_rst), .Q(n3348), .QN() );
  DFFR_X1 reg_b_reg_30_ ( .D(n1297), .CK(i_clk), .RN(i_rst), .Q(reg_b[30]), 
        .QN(n701) );
  DFFR_X1 sdata_reg_31_ ( .D(n1296), .CK(i_clk), .RN(i_rst), .Q(sdata[31]), 
        .QN(n2814) );
  DFFR_X1 state_reg_5_ ( .D(n1229), .CK(i_clk), .RN(i_rst), .Q(state[5]), 
        .QN() );
  DFFR_X1 state_reg_4_ ( .D(n1192), .CK(i_clk), .RN(i_rst), .Q(state[4]), .QN(
        n2806) );
  DFFS_X1 state_reg_0_ ( .D(n1191), .CK(i_clk), .SN(i_rst), .Q(state[0]), .QN(
        n2807) );
  DFFR_X1 state_reg_1_ ( .D(n1228), .CK(i_clk), .RN(i_rst), .Q(state[1]), .QN(
        n2799) );
  DFFR_X1 state_reg_2_ ( .D(n1226), .CK(i_clk), .RN(i_rst), .Q(state[2]), .QN(
        n2855) );
  DFFR_X1 state_reg_3_ ( .D(n1225), .CK(i_clk), .RN(i_rst), .Q(state[3]), .QN(
        n2853) );
  DFFR_X1 o_quotient_reg_31_ ( .D(n1193), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[31]), .QN() );
  DFFR_X1 o_quotient_reg_30_ ( .D(n1194), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[30]), .QN() );
  DFFR_X1 o_quotient_reg_29_ ( .D(n1195), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[29]), .QN() );
  DFFR_X1 o_quotient_reg_28_ ( .D(n1196), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[28]), .QN() );
  DFFR_X1 o_quotient_reg_27_ ( .D(n1197), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[27]), .QN() );
  DFFR_X1 o_quotient_reg_26_ ( .D(n1198), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[26]), .QN() );
  DFFR_X1 o_quotient_reg_25_ ( .D(n1199), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[25]), .QN() );
  DFFR_X1 o_quotient_reg_24_ ( .D(n1200), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[24]), .QN() );
  DFFR_X1 o_quotient_reg_23_ ( .D(n1201), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[23]), .QN() );
  DFFR_X1 o_quotient_reg_22_ ( .D(n1202), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[22]), .QN() );
  DFFR_X1 o_quotient_reg_21_ ( .D(n1203), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[21]), .QN() );
  DFFR_X1 o_quotient_reg_20_ ( .D(n1204), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[20]), .QN() );
  DFFR_X1 o_quotient_reg_19_ ( .D(n1205), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[19]), .QN() );
  DFFR_X1 o_quotient_reg_18_ ( .D(n1206), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[18]), .QN() );
  DFFR_X1 o_quotient_reg_17_ ( .D(n1207), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[17]), .QN() );
  DFFR_X1 o_quotient_reg_16_ ( .D(n1208), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[16]), .QN() );
  DFFR_X1 o_quotient_reg_15_ ( .D(n1209), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[15]), .QN() );
  DFFR_X1 o_quotient_reg_14_ ( .D(n1210), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[14]), .QN() );
  DFFR_X1 o_quotient_reg_13_ ( .D(n1211), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[13]), .QN() );
  DFFR_X1 o_quotient_reg_12_ ( .D(n1212), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[12]), .QN() );
  DFFR_X1 o_quotient_reg_11_ ( .D(n1213), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[11]), .QN() );
  DFFR_X1 o_quotient_reg_10_ ( .D(n1214), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[10]), .QN() );
  DFFR_X1 o_quotient_reg_9_ ( .D(n1215), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[9]), .QN() );
  DFFR_X1 o_quotient_reg_8_ ( .D(n1216), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[8]), .QN() );
  DFFR_X1 o_quotient_reg_7_ ( .D(n1217), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[7]), .QN() );
  DFFR_X1 o_quotient_reg_6_ ( .D(n1218), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[6]), .QN() );
  DFFR_X1 o_quotient_reg_5_ ( .D(n1219), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[5]), .QN() );
  DFFR_X1 o_quotient_reg_4_ ( .D(n1220), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[4]), .QN() );
  DFFR_X1 o_quotient_reg_3_ ( .D(n1221), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[3]), .QN() );
  DFFR_X1 o_quotient_reg_2_ ( .D(n1222), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[2]), .QN() );
  DFFR_X1 o_quotient_reg_1_ ( .D(n1223), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[1]), .QN() );
  DFFR_X1 o_quotient_reg_0_ ( .D(n1224), .CK(i_clk), .RN(i_rst), .Q(
        o_quotient[0]), .QN() );
  SDFFR_X1 state_reg_reg_1_ ( .D(1'b1), .SI(n977), .SE(n941), .CK(i_clk), .RN(
        i_rst), .Q(state_reg_1_0), .QN() );
  DFFR_X1 state_reg_reg_0_ ( .D(n1293), .CK(i_clk), .RN(i_rst), .Q(n3347), 
        .QN(n941) );
  DFFR_X1 ready_reg ( .D(n1230), .CK(i_clk), .RN(i_rst), .Q(ready), .QN(n2817)
         );
  DFFR_X1 o_remainder_reg_31_ ( .D(n1231), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[31]), .QN() );
  DFFR_X1 o_remainder_reg_30_ ( .D(n1232), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[30]), .QN() );
  DFFR_X1 o_remainder_reg_29_ ( .D(n1233), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[29]), .QN() );
  DFFR_X1 o_remainder_reg_28_ ( .D(n1234), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[28]), .QN() );
  DFFR_X1 o_remainder_reg_27_ ( .D(n1235), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[27]), .QN() );
  DFFR_X1 o_remainder_reg_26_ ( .D(n1236), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[26]), .QN() );
  DFFR_X1 o_remainder_reg_25_ ( .D(n1237), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[25]), .QN() );
  DFFR_X1 o_remainder_reg_24_ ( .D(n1238), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[24]), .QN() );
  DFFR_X1 o_remainder_reg_23_ ( .D(n1239), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[23]), .QN() );
  DFFR_X1 o_remainder_reg_22_ ( .D(n1240), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[22]), .QN() );
  DFFR_X1 o_remainder_reg_21_ ( .D(n1241), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[21]), .QN() );
  DFFR_X1 o_remainder_reg_20_ ( .D(n1242), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[20]), .QN() );
  DFFR_X1 o_remainder_reg_19_ ( .D(n1243), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[19]), .QN() );
  DFFR_X1 o_remainder_reg_18_ ( .D(n1244), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[18]), .QN() );
  DFFR_X1 o_remainder_reg_17_ ( .D(n1245), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[17]), .QN() );
  DFFR_X1 o_remainder_reg_16_ ( .D(n1246), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[16]), .QN() );
  DFFR_X1 o_remainder_reg_15_ ( .D(n1247), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[15]), .QN() );
  DFFR_X1 o_remainder_reg_14_ ( .D(n1248), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[14]), .QN() );
  DFFR_X1 o_remainder_reg_13_ ( .D(n1249), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[13]), .QN() );
  DFFR_X1 o_remainder_reg_12_ ( .D(n1250), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[12]), .QN() );
  DFFR_X1 o_remainder_reg_11_ ( .D(n1251), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[11]), .QN() );
  DFFR_X1 o_remainder_reg_10_ ( .D(n1252), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[10]), .QN() );
  DFFR_X1 o_remainder_reg_9_ ( .D(n1253), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[9]), .QN() );
  DFFR_X1 o_remainder_reg_8_ ( .D(n1254), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[8]), .QN() );
  DFFR_X1 o_remainder_reg_7_ ( .D(n1255), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[7]), .QN() );
  DFFR_X1 o_remainder_reg_6_ ( .D(n1256), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[6]), .QN() );
  DFFR_X1 o_remainder_reg_5_ ( .D(n1257), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[5]), .QN() );
  DFFR_X1 o_remainder_reg_4_ ( .D(n1258), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[4]), .QN() );
  DFFR_X1 o_remainder_reg_3_ ( .D(n1259), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[3]), .QN() );
  DFFR_X1 o_remainder_reg_2_ ( .D(n1260), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[2]), .QN() );
  DFFR_X1 o_remainder_reg_1_ ( .D(n1261), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[1]), .QN() );
  DFFR_X1 o_remainder_reg_0_ ( .D(n1262), .CK(i_clk), .RN(i_rst), .Q(
        o_remainder[0]), .QN() );
  DFFR_X1 DD_sign_reg ( .D(n1227), .CK(i_clk), .RN(i_rst), .Q(n3272), .QN(
        n2854) );
  DFFR_X1 ct_reg_5_ ( .D(n3358), .CK(i_clk), .RN(i_rst), .Q(ct[5]), .QN(n934)
         );
  DFFR_X1 sdata_reg_0_ ( .D(n1186), .CK(i_clk), .RN(i_rst), .Q(sdata[0]), .QN(
        n2825) );
  DFFR_X1 shifted_reg_0_ ( .D(n1190), .CK(i_clk), .RN(i_rst), .Q(), .QN(n3346)
         );
  DFFR_X1 shifted_reg_1_ ( .D(n1189), .CK(i_clk), .RN(i_rst), .Q(), .QN(n3345)
         );
  DFFR_X1 shifted_reg_2_ ( .D(n1188), .CK(i_clk), .RN(i_rst), .Q(), .QN(n3344)
         );
  DFFR_X1 shifted_reg_3_ ( .D(n1187), .CK(i_clk), .RN(i_rst), .Q(), .QN(n3343)
         );
  DFFR_X1 PR_reg_1_ ( .D(n3354), .CK(i_clk), .RN(i_rst), .Q(n3342), .QN() );
  DFFR_X1 sdata_reg_1_ ( .D(n1185), .CK(i_clk), .RN(i_rst), .Q(sdata[1]), .QN(
        n2826) );
  DFFR_X1 DR_reg_1_ ( .D(n1154), .CK(i_clk), .RN(i_rst), .Q(n3341), .QN() );
  DFFR_X1 PR_reg_2_ ( .D(n3353), .CK(i_clk), .RN(i_rst), .Q(n3340), .QN() );
  DFFR_X1 sdata_reg_2_ ( .D(n1184), .CK(i_clk), .RN(i_rst), .Q(sdata[2]), .QN(
        n2827) );
  DFFR_X1 DR_reg_2_ ( .D(n1153), .CK(i_clk), .RN(i_rst), .Q(n3339), .QN() );
  DFFR_X1 PR_reg_3_ ( .D(n3351), .CK(i_clk), .RN(i_rst), .Q(n3338), .QN() );
  DFFR_X1 sdata_reg_3_ ( .D(n1183), .CK(i_clk), .RN(i_rst), .Q(sdata[3]), .QN(
        n2828) );
  DFFR_X1 DR_reg_3_ ( .D(n1152), .CK(i_clk), .RN(i_rst), .Q(n3337), .QN() );
  DFFR_X1 PR_reg_4_ ( .D(n3350), .CK(i_clk), .RN(i_rst), .Q(n3336), .QN() );
  DFFR_X1 sdata_reg_4_ ( .D(n1182), .CK(i_clk), .RN(i_rst), .Q(sdata[4]), .QN(
        n2829) );
  DFFR_X1 DR_reg_4_ ( .D(n1151), .CK(i_clk), .RN(i_rst), .Q(n3335), .QN() );
  DFFR_X1 PR_reg_5_ ( .D(n3349), .CK(i_clk), .RN(i_rst), .Q(n3334), .QN() );
  DFFR_X1 sdata_reg_5_ ( .D(n1181), .CK(i_clk), .RN(i_rst), .Q(sdata[5]), .QN(
        n2830) );
  DFFR_X1 DR_reg_5_ ( .D(n1150), .CK(i_clk), .RN(i_rst), .Q(n3333), .QN() );
  DFFR_X1 PR_reg_6_ ( .D(n862), .CK(i_clk), .RN(i_rst), .Q(n3285), .QN(n2787)
         );
  DFFR_X1 sdata_reg_6_ ( .D(n1180), .CK(i_clk), .RN(i_rst), .Q(sdata[6]), .QN(
        n2831) );
  DFFR_X1 DR_reg_6_ ( .D(n1149), .CK(i_clk), .RN(i_rst), .Q(n3332), .QN() );
  DFFR_X1 PR_reg_7_ ( .D(n861), .CK(i_clk), .RN(i_rst), .Q(n3284), .QN(n2848)
         );
  DFFR_X1 sdata_reg_7_ ( .D(n1179), .CK(i_clk), .RN(i_rst), .Q(sdata[7]), .QN(
        n2832) );
  DFFR_X1 DR_reg_7_ ( .D(n1148), .CK(i_clk), .RN(i_rst), .Q(n3331), .QN() );
  DFFR_X1 PR_reg_8_ ( .D(n860), .CK(i_clk), .RN(i_rst), .Q(n3283), .QN(n2801)
         );
  DFFR_X1 sdata_reg_8_ ( .D(n1178), .CK(i_clk), .RN(i_rst), .Q(sdata[8]), .QN(
        n2833) );
  DFFR_X1 DR_reg_8_ ( .D(n1147), .CK(i_clk), .RN(i_rst), .Q(n3330), .QN() );
  DFFR_X1 PR_reg_9_ ( .D(n859), .CK(i_clk), .RN(i_rst), .Q(n3282), .QN(n2794)
         );
  DFFR_X1 sdata_reg_9_ ( .D(n1177), .CK(i_clk), .RN(i_rst), .Q(sdata[9]), .QN(
        n2834) );
  DFFR_X1 DR_reg_9_ ( .D(n1146), .CK(i_clk), .RN(i_rst), .Q(n3329), .QN() );
  DFFR_X1 PR_reg_10_ ( .D(n858), .CK(i_clk), .RN(i_rst), .Q(n3289), .QN(n2792)
         );
  DFFR_X1 sdata_reg_10_ ( .D(n1176), .CK(i_clk), .RN(i_rst), .Q(sdata[10]), 
        .QN(n2835) );
  DFFR_X1 DR_reg_10_ ( .D(n1145), .CK(i_clk), .RN(i_rst), .Q(n3328), .QN() );
  DFFR_X1 PR_reg_11_ ( .D(n857), .CK(i_clk), .RN(i_rst), .Q(n3288), .QN(n2847)
         );
  DFFR_X1 sdata_reg_11_ ( .D(n1175), .CK(i_clk), .RN(i_rst), .Q(sdata[11]), 
        .QN(n2836) );
  DFFR_X1 DR_reg_11_ ( .D(n1144), .CK(i_clk), .RN(i_rst), .Q(n3327), .QN() );
  DFFR_X1 PR_reg_12_ ( .D(n856), .CK(i_clk), .RN(i_rst), .Q(n3287), .QN(n2800)
         );
  DFFR_X1 sdata_reg_12_ ( .D(n1174), .CK(i_clk), .RN(i_rst), .Q(sdata[12]), 
        .QN(n2837) );
  DFFR_X1 DR_reg_12_ ( .D(n1143), .CK(i_clk), .RN(i_rst), .Q(n3326), .QN() );
  DFFR_X1 PR_reg_13_ ( .D(n855), .CK(i_clk), .RN(i_rst), .Q(n3286), .QN(n2793)
         );
  DFFR_X1 sdata_reg_13_ ( .D(n1173), .CK(i_clk), .RN(i_rst), .Q(sdata[13]), 
        .QN(n2838) );
  DFFR_X1 DR_reg_13_ ( .D(n1142), .CK(i_clk), .RN(i_rst), .Q(n3325), .QN() );
  DFFR_X1 PR_reg_14_ ( .D(n854), .CK(i_clk), .RN(i_rst), .Q(n3293), .QN(n2791)
         );
  DFFR_X1 sdata_reg_14_ ( .D(n1172), .CK(i_clk), .RN(i_rst), .Q(sdata[14]), 
        .QN(n2839) );
  DFFR_X1 DR_reg_14_ ( .D(n1141), .CK(i_clk), .RN(i_rst), .Q(n3324), .QN() );
  DFFR_X1 PR_reg_15_ ( .D(n853), .CK(i_clk), .RN(i_rst), .Q(n3292), .QN(n2852)
         );
  DFFR_X1 sdata_reg_15_ ( .D(n1171), .CK(i_clk), .RN(i_rst), .Q(sdata[15]), 
        .QN(n2840) );
  DFFR_X1 DR_reg_15_ ( .D(n1140), .CK(i_clk), .RN(i_rst), .Q(n3323), .QN() );
  DFFR_X1 PR_reg_16_ ( .D(n852), .CK(i_clk), .RN(i_rst), .Q(n3291), .QN(n2805)
         );
  DFFR_X1 sdata_reg_16_ ( .D(n1170), .CK(i_clk), .RN(i_rst), .Q(sdata[16]), 
        .QN(n2841) );
  DFFR_X1 DR_reg_16_ ( .D(n1139), .CK(i_clk), .RN(i_rst), .Q(n3322), .QN() );
  DFFR_X1 PR_reg_17_ ( .D(n851), .CK(i_clk), .RN(i_rst), .Q(n3290), .QN(n2798)
         );
  DFFR_X1 sdata_reg_17_ ( .D(n1169), .CK(i_clk), .RN(i_rst), .Q(sdata[17]), 
        .QN(n2842) );
  DFFR_X1 DR_reg_17_ ( .D(n1138), .CK(i_clk), .RN(i_rst), .Q(n3321), .QN() );
  DFFR_X1 PR_reg_18_ ( .D(n850), .CK(i_clk), .RN(i_rst), .Q(n3297), .QN(n2858)
         );
  DFFR_X1 sdata_reg_18_ ( .D(n1168), .CK(i_clk), .RN(i_rst), .Q(sdata[18]), 
        .QN(n2843) );
  DFFR_X1 DR_reg_18_ ( .D(n1137), .CK(i_clk), .RN(i_rst), .Q(n3320), .QN() );
  DFFR_X1 PR_reg_19_ ( .D(n849), .CK(i_clk), .RN(i_rst), .Q(n3296), .QN(n2851)
         );
  DFFR_X1 sdata_reg_19_ ( .D(n1167), .CK(i_clk), .RN(i_rst), .Q(sdata[19]), 
        .QN(n2844) );
  DFFR_X1 DR_reg_19_ ( .D(n1136), .CK(i_clk), .RN(i_rst), .Q(n3319), .QN() );
  DFFR_X1 PR_reg_20_ ( .D(n848), .CK(i_clk), .RN(i_rst), .Q(n3295), .QN(n2804)
         );
  DFFR_X1 sdata_reg_20_ ( .D(n1166), .CK(i_clk), .RN(i_rst), .Q(sdata[20]), 
        .QN(n2845) );
  DFFR_X1 DR_reg_20_ ( .D(n1135), .CK(i_clk), .RN(i_rst), .Q(n3318), .QN() );
  DFFR_X1 PR_reg_21_ ( .D(n847), .CK(i_clk), .RN(i_rst), .Q(n3294), .QN(n2797)
         );
  DFFR_X1 sdata_reg_21_ ( .D(n1165), .CK(i_clk), .RN(i_rst), .Q(sdata[21]), 
        .QN(n2846) );
  DFFR_X1 DR_reg_21_ ( .D(n1134), .CK(i_clk), .RN(i_rst), .Q(n3317), .QN() );
  DFFR_X1 PR_reg_22_ ( .D(n846), .CK(i_clk), .RN(i_rst), .Q(n3276), .QN(n2850)
         );
  DFFR_X1 sdata_reg_22_ ( .D(n1164), .CK(i_clk), .RN(i_rst), .Q(sdata[22]), 
        .QN(n2818) );
  DFFR_X1 DR_reg_22_ ( .D(n1133), .CK(i_clk), .RN(i_rst), .Q(n3316), .QN() );
  DFFR_X1 PR_reg_23_ ( .D(n845), .CK(i_clk), .RN(i_rst), .Q(n3275), .QN(n2803)
         );
  DFFR_X1 sdata_reg_23_ ( .D(n1163), .CK(i_clk), .RN(i_rst), .Q(sdata[23]), 
        .QN(n2819) );
  DFFR_X1 DR_reg_23_ ( .D(n1132), .CK(i_clk), .RN(i_rst), .Q(n3315), .QN() );
  DFFR_X1 PR_reg_24_ ( .D(n844), .CK(i_clk), .RN(i_rst), .Q(n3274), .QN(n2796)
         );
  DFFR_X1 sdata_reg_24_ ( .D(n1162), .CK(i_clk), .RN(i_rst), .Q(sdata[24]), 
        .QN(n2820) );
  DFFR_X1 DR_reg_24_ ( .D(n1131), .CK(i_clk), .RN(i_rst), .Q(n3314), .QN() );
  DFFR_X1 PR_reg_25_ ( .D(n843), .CK(i_clk), .RN(i_rst), .Q(n3273), .QN(n2790)
         );
  DFFR_X1 sdata_reg_25_ ( .D(n1161), .CK(i_clk), .RN(i_rst), .Q(sdata[25]), 
        .QN(n2824) );
  DFFR_X1 DR_reg_25_ ( .D(n1130), .CK(i_clk), .RN(i_rst), .Q(n3313), .QN() );
  DFFR_X1 PR_reg_26_ ( .D(n842), .CK(i_clk), .RN(i_rst), .Q(n3280), .QN(n2849)
         );
  DFFR_X1 sdata_reg_26_ ( .D(n1160), .CK(i_clk), .RN(i_rst), .Q(sdata[26]), 
        .QN(n2815) );
  DFFR_X1 DR_reg_26_ ( .D(n1129), .CK(i_clk), .RN(i_rst), .Q(n3312), .QN() );
  DFFR_X1 PR_reg_27_ ( .D(n841), .CK(i_clk), .RN(i_rst), .Q(n3279), .QN(n2802)
         );
  DFFR_X1 sdata_reg_27_ ( .D(n1159), .CK(i_clk), .RN(i_rst), .Q(sdata[27]), 
        .QN(n2821) );
  DFFR_X1 DR_reg_27_ ( .D(n1128), .CK(i_clk), .RN(i_rst), .Q(n3311), .QN() );
  DFFR_X1 PR_reg_28_ ( .D(n840), .CK(i_clk), .RN(i_rst), .Q(n3278), .QN(n2795)
         );
  DFFR_X1 sdata_reg_28_ ( .D(n1158), .CK(i_clk), .RN(i_rst), .Q(sdata[28]), 
        .QN(n2822) );
  DFFR_X1 DR_reg_28_ ( .D(n1127), .CK(i_clk), .RN(i_rst), .Q(n3310), .QN() );
  DFFR_X1 PR_reg_29_ ( .D(n839), .CK(i_clk), .RN(i_rst), .Q(n3277), .QN(n2789)
         );
  DFFR_X1 sdata_reg_29_ ( .D(n1157), .CK(i_clk), .RN(i_rst), .Q(sdata[29]), 
        .QN(n2823) );
  DFFR_X1 DR_reg_29_ ( .D(n1126), .CK(i_clk), .RN(i_rst), .Q(n3309), .QN() );
  DFFR_X1 PR_reg_30_ ( .D(n838), .CK(i_clk), .RN(i_rst), .Q(n3281), .QN(n2788)
         );
  DFFR_X1 sdata_reg_30_ ( .D(n1156), .CK(i_clk), .RN(i_rst), .Q(sdata[30]), 
        .QN(n2816) );
  DFFR_X1 DR_reg_30_ ( .D(n1125), .CK(i_clk), .RN(i_rst), .Q(n3308), .QN() );
  DFFR_X1 PR_reg_31_ ( .D(n3352), .CK(i_clk), .RN(i_rst), .Q(n2856), .QN(n3307) );
  DFFR_X1 DR_reg_0_ ( .D(n1155), .CK(i_clk), .RN(i_rst), .Q(n3306), .QN() );
  DFFR_X1 ct_1_en_reg ( .D(n1113), .CK(i_clk), .RN(i_rst), .Q(n3298), .QN() );
  DFFR_X1 ct_1_en_1_reg ( .D(n1864), .CK(i_clk), .RN(i_rst), .Q(), .QN(n3305)
         );
  DFFR_X1 ct_1_reg_5_ ( .D(n1106), .CK(i_clk), .RN(i_rst), .Q(ct_1[5]), .QN(
        n944) );
  DFFR_X1 ct_1_reg_4_ ( .D(n1107), .CK(i_clk), .RN(i_rst), .Q(ct_1[4]), .QN(
        n945) );
  DFFR_X1 ct_1_reg_3_ ( .D(n1108), .CK(i_clk), .RN(i_rst), .Q(ct_1[3]), .QN(
        n946) );
  DFFR_X1 ct_1_reg_2_ ( .D(n1109), .CK(i_clk), .RN(i_rst), .Q(ct_1[2]), .QN(
        n947) );
  DFFR_X1 ct_1_reg_1_ ( .D(n1110), .CK(i_clk), .RN(i_rst), .Q(ct_1[1]), .QN(
        n948) );
  DFFR_X1 ct_1_reg_0_ ( .D(n1111), .CK(i_clk), .RN(i_rst), .Q(ct_1[0]), .QN(
        n949) );
  DFFR_X1 shifted_1_reg_3_ ( .D(n2786), .CK(i_clk), .RN(i_rst), .Q(), .QN(
        n3304) );
  DFFR_X1 shifted_1_reg_2_ ( .D(n2785), .CK(i_clk), .RN(i_rst), .Q(), .QN(
        n3303) );
  DFFR_X1 shifted_1_reg_1_ ( .D(n2784), .CK(i_clk), .RN(i_rst), .Q(), .QN(
        n3302) );
  DFFR_X1 shifted_1_reg_0_ ( .D(n2783), .CK(i_clk), .RN(i_rst), .Q(), .QN(
        n3301) );
  DFFR_X1 ct_reg_4_ ( .D(n3356), .CK(i_clk), .RN(i_rst), .Q(ct[4]), .QN(n935)
         );
  DFFR_X1 ct_reg_3_ ( .D(n3357), .CK(i_clk), .RN(i_rst), .Q(ct[3]), .QN(n936)
         );
  DFFR_X1 ct_reg_2_ ( .D(n3359), .CK(i_clk), .RN(i_rst), .Q(ct[2]), .QN(n937)
         );
  DFFR_X1 ct_reg_1_ ( .D(n3360), .CK(i_clk), .RN(i_rst), .Q(ct[1]), .QN(n938)
         );
  DFFR_X1 ct_reg_0_ ( .D(n3361), .CK(i_clk), .RN(i_rst), .Q(ct[0]), .QN(n939)
         );
  DFFR_X1 DR_reg_31_ ( .D(n1124), .CK(i_clk), .RN(i_rst), .Q(n3299), .QN() );
  DFFR_X1 reg_carry_reg ( .D(n1043), .CK(i_clk), .RN(i_rst), .Q(reg_carry), 
        .QN(n940) );
  DFFR_X1 q_reg_30_ ( .D(n1044), .CK(i_clk), .RN(i_rst), .Q(q[30]), .QN() );
  DFFR_X1 q_reg_29_ ( .D(n1045), .CK(i_clk), .RN(i_rst), .Q(q[29]), .QN() );
  DFFR_X1 q_reg_28_ ( .D(n1046), .CK(i_clk), .RN(i_rst), .Q(q[28]), .QN() );
  DFFR_X1 q_reg_27_ ( .D(n1047), .CK(i_clk), .RN(i_rst), .Q(q[27]), .QN() );
  DFFR_X1 q_reg_26_ ( .D(n1048), .CK(i_clk), .RN(i_rst), .Q(q[26]), .QN() );
  DFFR_X1 q_reg_25_ ( .D(n1049), .CK(i_clk), .RN(i_rst), .Q(q[25]), .QN() );
  DFFR_X1 q_reg_24_ ( .D(n1050), .CK(i_clk), .RN(i_rst), .Q(q[24]), .QN() );
  DFFR_X1 q_reg_23_ ( .D(n1051), .CK(i_clk), .RN(i_rst), .Q(q[23]), .QN() );
  DFFR_X1 q_reg_22_ ( .D(n1052), .CK(i_clk), .RN(i_rst), .Q(q[22]), .QN() );
  DFFR_X1 q_reg_21_ ( .D(n1053), .CK(i_clk), .RN(i_rst), .Q(q[21]), .QN() );
  DFFR_X1 q_reg_20_ ( .D(n1054), .CK(i_clk), .RN(i_rst), .Q(q[20]), .QN() );
  DFFR_X1 q_reg_19_ ( .D(n1055), .CK(i_clk), .RN(i_rst), .Q(q[19]), .QN() );
  DFFR_X1 q_reg_18_ ( .D(n1056), .CK(i_clk), .RN(i_rst), .Q(q[18]), .QN() );
  DFFR_X1 q_reg_17_ ( .D(n1057), .CK(i_clk), .RN(i_rst), .Q(q[17]), .QN() );
  DFFR_X1 q_reg_16_ ( .D(n1058), .CK(i_clk), .RN(i_rst), .Q(q[16]), .QN() );
  DFFR_X1 q_reg_15_ ( .D(n1059), .CK(i_clk), .RN(i_rst), .Q(q[15]), .QN() );
  DFFR_X1 q_reg_14_ ( .D(n1060), .CK(i_clk), .RN(i_rst), .Q(q[14]), .QN() );
  DFFR_X1 q_reg_13_ ( .D(n1061), .CK(i_clk), .RN(i_rst), .Q(q[13]), .QN() );
  DFFR_X1 q_reg_12_ ( .D(n1062), .CK(i_clk), .RN(i_rst), .Q(q[12]), .QN() );
  DFFR_X1 q_reg_11_ ( .D(n1063), .CK(i_clk), .RN(i_rst), .Q(q[11]), .QN() );
  DFFR_X1 q_reg_10_ ( .D(n1064), .CK(i_clk), .RN(i_rst), .Q(q[10]), .QN() );
  DFFR_X1 q_reg_9_ ( .D(n1065), .CK(i_clk), .RN(i_rst), .Q(q[9]), .QN() );
  DFFR_X1 q_reg_8_ ( .D(n1066), .CK(i_clk), .RN(i_rst), .Q(q[8]), .QN() );
  DFFR_X1 q_reg_7_ ( .D(n1067), .CK(i_clk), .RN(i_rst), .Q(q[7]), .QN() );
  DFFR_X1 q_reg_6_ ( .D(n1068), .CK(i_clk), .RN(i_rst), .Q(q[6]), .QN() );
  DFFR_X1 q_reg_5_ ( .D(n1069), .CK(i_clk), .RN(i_rst), .Q(q[5]), .QN() );
  DFFR_X1 q_reg_4_ ( .D(n1070), .CK(i_clk), .RN(i_rst), .Q(q[4]), .QN() );
  DFFR_X1 q_reg_3_ ( .D(n1071), .CK(i_clk), .RN(i_rst), .Q(q[3]), .QN() );
  DFFR_X1 q_reg_2_ ( .D(n1072), .CK(i_clk), .RN(i_rst), .Q(q[2]), .QN() );
  DFFR_X1 q_reg_1_ ( .D(n1073), .CK(i_clk), .RN(i_rst), .Q(q[1]), .QN() );
  DFFR_X1 q_reg_0_ ( .D(n1074), .CK(i_clk), .RN(i_rst), .Q(q[0]), .QN() );
  DFFR_X1 nq_reg_30_ ( .D(n1075), .CK(i_clk), .RN(i_rst), .Q(nq[30]), .QN() );
  DFFR_X1 nq_reg_29_ ( .D(n1076), .CK(i_clk), .RN(i_rst), .Q(nq[29]), .QN() );
  DFFR_X1 nq_reg_28_ ( .D(n1077), .CK(i_clk), .RN(i_rst), .Q(nq[28]), .QN() );
  DFFR_X1 nq_reg_27_ ( .D(n1078), .CK(i_clk), .RN(i_rst), .Q(nq[27]), .QN() );
  DFFR_X1 nq_reg_26_ ( .D(n1079), .CK(i_clk), .RN(i_rst), .Q(nq[26]), .QN() );
  DFFR_X1 nq_reg_25_ ( .D(n1080), .CK(i_clk), .RN(i_rst), .Q(nq[25]), .QN() );
  DFFR_X1 nq_reg_24_ ( .D(n1081), .CK(i_clk), .RN(i_rst), .Q(nq[24]), .QN() );
  DFFR_X1 nq_reg_23_ ( .D(n1082), .CK(i_clk), .RN(i_rst), .Q(nq[23]), .QN() );
  DFFR_X1 nq_reg_22_ ( .D(n1083), .CK(i_clk), .RN(i_rst), .Q(nq[22]), .QN() );
  DFFR_X1 nq_reg_21_ ( .D(n1084), .CK(i_clk), .RN(i_rst), .Q(nq[21]), .QN() );
  DFFR_X1 nq_reg_20_ ( .D(n1085), .CK(i_clk), .RN(i_rst), .Q(nq[20]), .QN() );
  DFFR_X1 nq_reg_19_ ( .D(n1086), .CK(i_clk), .RN(i_rst), .Q(nq[19]), .QN() );
  DFFR_X1 nq_reg_18_ ( .D(n1087), .CK(i_clk), .RN(i_rst), .Q(nq[18]), .QN() );
  DFFR_X1 nq_reg_17_ ( .D(n1088), .CK(i_clk), .RN(i_rst), .Q(nq[17]), .QN() );
  DFFR_X1 nq_reg_16_ ( .D(n1089), .CK(i_clk), .RN(i_rst), .Q(nq[16]), .QN() );
  DFFR_X1 nq_reg_15_ ( .D(n1090), .CK(i_clk), .RN(i_rst), .Q(nq[15]), .QN() );
  DFFR_X1 nq_reg_14_ ( .D(n1091), .CK(i_clk), .RN(i_rst), .Q(nq[14]), .QN() );
  DFFR_X1 nq_reg_13_ ( .D(n1092), .CK(i_clk), .RN(i_rst), .Q(nq[13]), .QN() );
  DFFR_X1 nq_reg_12_ ( .D(n1093), .CK(i_clk), .RN(i_rst), .Q(nq[12]), .QN() );
  DFFR_X1 nq_reg_11_ ( .D(n1094), .CK(i_clk), .RN(i_rst), .Q(nq[11]), .QN() );
  DFFR_X1 nq_reg_10_ ( .D(n1095), .CK(i_clk), .RN(i_rst), .Q(nq[10]), .QN() );
  DFFR_X1 nq_reg_9_ ( .D(n1096), .CK(i_clk), .RN(i_rst), .Q(nq[9]), .QN() );
  DFFR_X1 nq_reg_8_ ( .D(n1097), .CK(i_clk), .RN(i_rst), .Q(nq[8]), .QN() );
  DFFR_X1 nq_reg_7_ ( .D(n1098), .CK(i_clk), .RN(i_rst), .Q(nq[7]), .QN() );
  DFFR_X1 nq_reg_6_ ( .D(n1099), .CK(i_clk), .RN(i_rst), .Q(nq[6]), .QN() );
  DFFR_X1 nq_reg_5_ ( .D(n1100), .CK(i_clk), .RN(i_rst), .Q(nq[5]), .QN() );
  DFFR_X1 nq_reg_4_ ( .D(n1101), .CK(i_clk), .RN(i_rst), .Q(nq[4]), .QN() );
  DFFR_X1 nq_reg_3_ ( .D(n1102), .CK(i_clk), .RN(i_rst), .Q(nq[3]), .QN() );
  DFFR_X1 nq_reg_2_ ( .D(n1103), .CK(i_clk), .RN(i_rst), .Q(nq[2]), .QN() );
  DFFR_X1 nq_reg_1_ ( .D(n1104), .CK(i_clk), .RN(i_rst), .Q(nq[1]), .QN() );
  DFFR_X1 nq_reg_0_ ( .D(n1105), .CK(i_clk), .RN(i_rst), .Q(nq[0]), .QN() );
  DFFR_X1 reg_a_reg_1_ ( .D(n1041), .CK(i_clk), .RN(i_rst), .Q(reg_a[1]), .QN(
        n1772) );
  DFFR_X1 reg_a_reg_2_ ( .D(n1040), .CK(i_clk), .RN(i_rst), .Q(reg_a[2]), .QN(
        n1771) );
  DFFR_X1 reg_a_reg_3_ ( .D(n1039), .CK(i_clk), .RN(i_rst), .Q(reg_a[3]), .QN(
        n1770) );
  DFFR_X1 reg_a_reg_4_ ( .D(n1038), .CK(i_clk), .RN(i_rst), .Q(reg_a[4]), .QN(
        n1769) );
  DFFR_X1 reg_a_reg_5_ ( .D(n1037), .CK(i_clk), .RN(i_rst), .Q(reg_a[5]), .QN(
        n802) );
  DFFR_X1 reg_a_reg_6_ ( .D(n1036), .CK(i_clk), .RN(i_rst), .Q(reg_a[6]), .QN(
        n803) );
  DFFR_X1 reg_a_reg_7_ ( .D(n1035), .CK(i_clk), .RN(i_rst), .Q(reg_a[7]), .QN(
        n804) );
  DFFR_X1 reg_a_reg_8_ ( .D(n1034), .CK(i_clk), .RN(i_rst), .Q(reg_a[8]), .QN(
        n805) );
  DFFR_X1 reg_a_reg_9_ ( .D(n1033), .CK(i_clk), .RN(i_rst), .Q(reg_a[9]), .QN(
        n806) );
  DFFR_X1 reg_a_reg_10_ ( .D(n1032), .CK(i_clk), .RN(i_rst), .Q(reg_a[10]), 
        .QN(n807) );
  DFFR_X1 reg_a_reg_11_ ( .D(n1031), .CK(i_clk), .RN(i_rst), .Q(reg_a[11]), 
        .QN(n808) );
  DFFR_X1 reg_a_reg_12_ ( .D(n1030), .CK(i_clk), .RN(i_rst), .Q(reg_a[12]), 
        .QN(n809) );
  DFFR_X1 reg_a_reg_13_ ( .D(n1029), .CK(i_clk), .RN(i_rst), .Q(reg_a[13]), 
        .QN(n810) );
  DFFR_X1 reg_a_reg_14_ ( .D(n1028), .CK(i_clk), .RN(i_rst), .Q(reg_a[14]), 
        .QN(n811) );
  DFFR_X1 reg_a_reg_15_ ( .D(n1027), .CK(i_clk), .RN(i_rst), .Q(reg_a[15]), 
        .QN(n812) );
  DFFR_X1 reg_a_reg_16_ ( .D(n1026), .CK(i_clk), .RN(i_rst), .Q(reg_a[16]), 
        .QN(n813) );
  DFFR_X1 reg_a_reg_17_ ( .D(n1025), .CK(i_clk), .RN(i_rst), .Q(reg_a[17]), 
        .QN(n814) );
  DFFR_X1 reg_a_reg_18_ ( .D(n1024), .CK(i_clk), .RN(i_rst), .Q(reg_a[18]), 
        .QN(n815) );
  DFFR_X1 reg_a_reg_19_ ( .D(n1023), .CK(i_clk), .RN(i_rst), .Q(reg_a[19]), 
        .QN(n816) );
  DFFR_X1 reg_a_reg_20_ ( .D(n1022), .CK(i_clk), .RN(i_rst), .Q(reg_a[20]), 
        .QN(n817) );
  DFFR_X1 reg_a_reg_21_ ( .D(n1021), .CK(i_clk), .RN(i_rst), .Q(reg_a[21]), 
        .QN(n818) );
  DFFR_X1 reg_a_reg_22_ ( .D(n1020), .CK(i_clk), .RN(i_rst), .Q(reg_a[22]), 
        .QN(n819) );
  DFFR_X1 reg_a_reg_23_ ( .D(n1019), .CK(i_clk), .RN(i_rst), .Q(reg_a[23]), 
        .QN(n820) );
  DFFR_X1 reg_a_reg_24_ ( .D(n1018), .CK(i_clk), .RN(i_rst), .Q(reg_a[24]), 
        .QN(n821) );
  DFFR_X1 reg_a_reg_25_ ( .D(n1017), .CK(i_clk), .RN(i_rst), .Q(reg_a[25]), 
        .QN(n822) );
  DFFR_X1 reg_a_reg_26_ ( .D(n1016), .CK(i_clk), .RN(i_rst), .Q(reg_a[26]), 
        .QN(n823) );
  DFFR_X1 reg_a_reg_27_ ( .D(n1015), .CK(i_clk), .RN(i_rst), .Q(reg_a[27]), 
        .QN(n824) );
  DFFR_X1 reg_a_reg_28_ ( .D(n1014), .CK(i_clk), .RN(i_rst), .Q(reg_a[28]), 
        .QN(n825) );
  DFFR_X1 reg_a_reg_29_ ( .D(n1013), .CK(i_clk), .RN(i_rst), .Q(reg_a[29]), 
        .QN(n826) );
  DFFR_X1 reg_a_reg_30_ ( .D(n1012), .CK(i_clk), .RN(i_rst), .Q(reg_a[30]), 
        .QN(n827) );
  DFFR_X1 reg_a_reg_0_ ( .D(n1042), .CK(i_clk), .RN(i_rst), .Q(reg_a[0]), .QN(
        n1773) );
  DFFR_X1 reg_a_reg_31_ ( .D(n1011), .CK(i_clk), .RN(i_rst), .Q(reg_a[31]), 
        .QN(n2857) );
  DFFR_X1 PR_1_reg_31_ ( .D(n979), .CK(i_clk), .RN(i_rst), .Q(PR_1[31]), .QN(
        n870) );
  DFFR_X1 PR_1_reg_0_ ( .D(n1010), .CK(i_clk), .RN(i_rst), .Q(PR_1[0]), .QN()
         );
  DFFR_X1 reg_b_reg_0_ ( .D(n1292), .CK(i_clk), .RN(i_rst), .Q(reg_b[0]), 
        .QN() );
  DFFR_X1 PR_1_reg_1_ ( .D(n1009), .CK(i_clk), .RN(i_rst), .Q(PR_1[1]), .QN()
         );
  DFFR_X1 reg_b_reg_1_ ( .D(n1291), .CK(i_clk), .RN(i_rst), .Q(reg_b[1]), 
        .QN() );
  DFFR_X1 PR_1_reg_2_ ( .D(n1008), .CK(i_clk), .RN(i_rst), .Q(PR_1[2]), .QN()
         );
  DFFR_X1 reg_b_reg_2_ ( .D(n1290), .CK(i_clk), .RN(i_rst), .Q(reg_b[2]), 
        .QN() );
  DFFR_X1 PR_1_reg_3_ ( .D(n1007), .CK(i_clk), .RN(i_rst), .Q(PR_1[3]), .QN()
         );
  DFFR_X1 reg_b_reg_3_ ( .D(n1289), .CK(i_clk), .RN(i_rst), .Q(reg_b[3]), 
        .QN() );
  DFFR_X1 PR_1_reg_4_ ( .D(n1006), .CK(i_clk), .RN(i_rst), .Q(PR_1[4]), .QN()
         );
  DFFR_X1 reg_b_reg_4_ ( .D(n1288), .CK(i_clk), .RN(i_rst), .Q(reg_b[4]), 
        .QN() );
  DFFR_X1 PR_1_reg_5_ ( .D(n1005), .CK(i_clk), .RN(i_rst), .Q(PR_1[5]), .QN()
         );
  DFFR_X1 reg_b_reg_5_ ( .D(n1287), .CK(i_clk), .RN(i_rst), .Q(reg_b[5]), 
        .QN() );
  DFFR_X1 PR_1_reg_6_ ( .D(n1004), .CK(i_clk), .RN(i_rst), .Q(PR_1[6]), .QN()
         );
  DFFR_X1 reg_b_reg_6_ ( .D(n1286), .CK(i_clk), .RN(i_rst), .Q(reg_b[6]), .QN(
        n708) );
  DFFR_X1 PR_1_reg_7_ ( .D(n1003), .CK(i_clk), .RN(i_rst), .Q(PR_1[7]), .QN()
         );
  DFFR_X1 reg_b_reg_7_ ( .D(n1285), .CK(i_clk), .RN(i_rst), .Q(reg_b[7]), .QN(
        n709) );
  DFFR_X1 PR_1_reg_8_ ( .D(n1002), .CK(i_clk), .RN(i_rst), .Q(PR_1[8]), .QN()
         );
  DFFR_X1 reg_b_reg_8_ ( .D(n1284), .CK(i_clk), .RN(i_rst), .Q(reg_b[8]), .QN(
        n710) );
  DFFR_X1 PR_1_reg_9_ ( .D(n1001), .CK(i_clk), .RN(i_rst), .Q(PR_1[9]), .QN()
         );
  DFFR_X1 reg_b_reg_9_ ( .D(n1283), .CK(i_clk), .RN(i_rst), .Q(reg_b[9]), .QN(
        n711) );
  DFFR_X1 PR_1_reg_10_ ( .D(n1000), .CK(i_clk), .RN(i_rst), .Q(PR_1[10]), 
        .QN() );
  DFFR_X1 reg_b_reg_10_ ( .D(n1282), .CK(i_clk), .RN(i_rst), .Q(reg_b[10]), 
        .QN(n712) );
  DFFR_X1 PR_1_reg_11_ ( .D(n999), .CK(i_clk), .RN(i_rst), .Q(PR_1[11]), .QN()
         );
  DFFR_X1 reg_b_reg_11_ ( .D(n1281), .CK(i_clk), .RN(i_rst), .Q(reg_b[11]), 
        .QN(n713) );
  DFFR_X1 PR_1_reg_12_ ( .D(n998), .CK(i_clk), .RN(i_rst), .Q(PR_1[12]), .QN()
         );
  DFFR_X1 reg_b_reg_12_ ( .D(n1280), .CK(i_clk), .RN(i_rst), .Q(reg_b[12]), 
        .QN(n714) );
  DFFR_X1 PR_1_reg_13_ ( .D(n997), .CK(i_clk), .RN(i_rst), .Q(PR_1[13]), .QN()
         );
  DFFR_X1 reg_b_reg_13_ ( .D(n1279), .CK(i_clk), .RN(i_rst), .Q(reg_b[13]), 
        .QN(n715) );
  DFFR_X1 PR_1_reg_14_ ( .D(n996), .CK(i_clk), .RN(i_rst), .Q(PR_1[14]), .QN()
         );
  DFFR_X1 reg_b_reg_14_ ( .D(n1278), .CK(i_clk), .RN(i_rst), .Q(reg_b[14]), 
        .QN(n716) );
  DFFR_X1 PR_1_reg_15_ ( .D(n995), .CK(i_clk), .RN(i_rst), .Q(PR_1[15]), .QN()
         );
  DFFR_X1 reg_b_reg_15_ ( .D(n1277), .CK(i_clk), .RN(i_rst), .Q(reg_b[15]), 
        .QN(n717) );
  DFFR_X1 PR_1_reg_16_ ( .D(n994), .CK(i_clk), .RN(i_rst), .Q(PR_1[16]), .QN()
         );
  DFFR_X1 reg_b_reg_16_ ( .D(n1276), .CK(i_clk), .RN(i_rst), .Q(reg_b[16]), 
        .QN(n718) );
  DFFR_X1 PR_1_reg_17_ ( .D(n993), .CK(i_clk), .RN(i_rst), .Q(PR_1[17]), .QN()
         );
  DFFR_X1 reg_b_reg_17_ ( .D(n1275), .CK(i_clk), .RN(i_rst), .Q(reg_b[17]), 
        .QN(n719) );
  DFFR_X1 PR_1_reg_18_ ( .D(n992), .CK(i_clk), .RN(i_rst), .Q(PR_1[18]), .QN()
         );
  DFFR_X1 reg_b_reg_18_ ( .D(n1274), .CK(i_clk), .RN(i_rst), .Q(reg_b[18]), 
        .QN(n720) );
  DFFR_X1 PR_1_reg_19_ ( .D(n991), .CK(i_clk), .RN(i_rst), .Q(PR_1[19]), .QN()
         );
  DFFR_X1 reg_b_reg_19_ ( .D(n1273), .CK(i_clk), .RN(i_rst), .Q(reg_b[19]), 
        .QN(n721) );
  DFFR_X1 PR_1_reg_20_ ( .D(n990), .CK(i_clk), .RN(i_rst), .Q(PR_1[20]), .QN()
         );
  DFFR_X1 reg_b_reg_20_ ( .D(n1272), .CK(i_clk), .RN(i_rst), .Q(reg_b[20]), 
        .QN(n722) );
  DFFR_X1 PR_1_reg_21_ ( .D(n989), .CK(i_clk), .RN(i_rst), .Q(PR_1[21]), .QN()
         );
  DFFR_X1 reg_b_reg_21_ ( .D(n1271), .CK(i_clk), .RN(i_rst), .Q(reg_b[21]), 
        .QN(n723) );
  DFFR_X1 PR_1_reg_22_ ( .D(n988), .CK(i_clk), .RN(i_rst), .Q(PR_1[22]), .QN()
         );
  DFFR_X1 reg_b_reg_22_ ( .D(n1270), .CK(i_clk), .RN(i_rst), .Q(reg_b[22]), 
        .QN(n724) );
  DFFR_X1 PR_1_reg_23_ ( .D(n987), .CK(i_clk), .RN(i_rst), .Q(PR_1[23]), .QN()
         );
  DFFR_X1 reg_b_reg_23_ ( .D(n1269), .CK(i_clk), .RN(i_rst), .Q(reg_b[23]), 
        .QN(n725) );
  DFFR_X1 PR_1_reg_24_ ( .D(n986), .CK(i_clk), .RN(i_rst), .Q(PR_1[24]), .QN()
         );
  DFFR_X1 reg_b_reg_24_ ( .D(n1268), .CK(i_clk), .RN(i_rst), .Q(reg_b[24]), 
        .QN(n726) );
  DFFR_X1 PR_1_reg_25_ ( .D(n985), .CK(i_clk), .RN(i_rst), .Q(PR_1[25]), .QN()
         );
  DFFR_X1 reg_b_reg_25_ ( .D(n1267), .CK(i_clk), .RN(i_rst), .Q(reg_b[25]), 
        .QN(n727) );
  DFFR_X1 PR_1_reg_26_ ( .D(n984), .CK(i_clk), .RN(i_rst), .Q(PR_1[26]), .QN()
         );
  DFFR_X1 reg_b_reg_26_ ( .D(n1266), .CK(i_clk), .RN(i_rst), .Q(reg_b[26]), 
        .QN(n728) );
  DFFR_X1 PR_1_reg_27_ ( .D(n983), .CK(i_clk), .RN(i_rst), .Q(PR_1[27]), .QN()
         );
  DFFR_X1 reg_b_reg_27_ ( .D(n1265), .CK(i_clk), .RN(i_rst), .Q(reg_b[27]), 
        .QN(n729) );
  DFFR_X1 PR_1_reg_28_ ( .D(n982), .CK(i_clk), .RN(i_rst), .Q(PR_1[28]), .QN()
         );
  DFFR_X1 reg_b_reg_28_ ( .D(n1264), .CK(i_clk), .RN(i_rst), .Q(reg_b[28]), 
        .QN(n730) );
  DFFR_X1 PR_1_reg_29_ ( .D(n981), .CK(i_clk), .RN(i_rst), .Q(PR_1[29]), .QN()
         );
  DFFR_X1 reg_b_reg_29_ ( .D(n1263), .CK(i_clk), .RN(i_rst), .Q(reg_b[29]), 
        .QN(n731) );
  DFFR_X1 PR_1_reg_30_ ( .D(n980), .CK(i_clk), .RN(i_rst), .Q(PR_1[30]), .QN()
         );
  DFFR_X1 reg_b_reg_31_ ( .D(n978), .CK(i_clk), .RN(i_rst), .Q(reg_b[31]), 
        .QN(n829) );
  OAI222_X1 U2114 ( .A1(nqp1[4]), .A2(n3135), .B1(1'b1), .B2(n2933), .C1(nq[4]), .C2(n3136), .ZN(n3153) );
  OR2_X1 U2115 ( .A1(n2984), .A2(n2926), .ZN(n2808) );
  OR2_X1 U2116 ( .A1(n3232), .A2(n2926), .ZN(n2809) );
  OR2_X1 U2117 ( .A1(n3112), .A2(n2925), .ZN(n2810) );
  OR3_X1 U2118 ( .A1(n2866), .A2(n2989), .A3(n2884), .ZN(n2811) );
  OR2_X1 U2119 ( .A1(n2982), .A2(n2984), .ZN(n2812) );
  OR2_X1 U2120 ( .A1(n2982), .A2(n2983), .ZN(n2813) );
  AND2_X2 U2121 ( .A1(n2988), .A2(n2938), .ZN(n2941) );
  AND2_X2 U2122 ( .A1(n2991), .A2(n2938), .ZN(n2942) );
  AND2_X2 U2123 ( .A1(n2990), .A2(n2938), .ZN(n2940) );
  NAND2_X2 U2124 ( .A1(n2986), .A2(n2938), .ZN(n2936) );
  INV_X1 U2125 ( .A(n2809), .ZN(n2859) );
  INV_X1 U2126 ( .A(n2810), .ZN(n2860) );
  INV_X1 U2127 ( .A(n2808), .ZN(n2861) );
  NOR2_X4 U2128 ( .A1(n2925), .A2(n3127), .ZN(n3137) );
  INV_X2 U2129 ( .A(n2947), .ZN(n2925) );
  NAND4_X2 U2130 ( .A1(n2995), .A2(n2875), .A3(n2943), .A4(n2881), .ZN(n2938)
         );
  INV_X2 U2131 ( .A(n2813), .ZN(n2862) );
  INV_X2 U2132 ( .A(n2812), .ZN(n2863) );
  INV_X2 U2133 ( .A(n2811), .ZN(n2864) );
  INV_X4 U2134 ( .A(n2997), .ZN(n2884) );
  NAND2_X4 U2135 ( .A1(n2876), .A2(n2880), .ZN(n2927) );
  NAND2_X2 U2136 ( .A1(n2990), .A2(n2998), .ZN(n2881) );
  OR2_X2 U2137 ( .A1(n3232), .A2(n2982), .ZN(n3135) );
  NAND2_X2 U2138 ( .A1(n2993), .A2(n2998), .ZN(n2985) );
  NOR2_X2 U2139 ( .A1(n3112), .A2(n2878), .ZN(n3080) );
  NAND2_X2 U2140 ( .A1(n3233), .A2(n3232), .ZN(n3136) );
  OR2_X2 U2141 ( .A1(n2875), .A2(n3068), .ZN(n2994) );
  NOR2_X2 U2142 ( .A1(n2878), .A2(n3127), .ZN(n3113) );
  NAND4_X2 U2143 ( .A1(n2986), .A2(n2998), .A3(i_start), .A4(n2817), .ZN(n2995) );
  NOR2_X4 U2144 ( .A1(n3129), .A2(n3130), .ZN(n2935) );
  INV_X2 U2145 ( .A(n2866), .ZN(n2880) );
  NOR2_X4 U2146 ( .A1(n941), .A2(state_reg_1_0), .ZN(n2866) );
  INV_X4 U2147 ( .A(state[5]), .ZN(n1988) );
  INV_X1 U2149 ( .A(n2865), .ZN(o_ready) );
  MUX2_X1 U2150 ( .A(n3334), .B(sdata_o[5]), .S(n2866), .Z(n3349) );
  MUX2_X1 U2151 ( .A(n3336), .B(sdata_o[4]), .S(n2866), .Z(n3350) );
  MUX2_X1 U2152 ( .A(n3338), .B(sdata_o[3]), .S(n2866), .Z(n3351) );
  MUX2_X1 U2153 ( .A(n2856), .B(sdata_o[31]), .S(n2866), .Z(n3352) );
  MUX2_X1 U2154 ( .A(n3340), .B(sdata_o[2]), .S(n2866), .Z(n3353) );
  MUX2_X1 U2155 ( .A(n3342), .B(sdata_o[1]), .S(n2866), .Z(n3354) );
  MUX2_X1 U2156 ( .A(n3348), .B(sdata_o[0]), .S(n2866), .Z(n3355) );
  INV_X1 U2157 ( .A(n2867), .ZN(n3356) );
  AOI22_X1 U2158 ( .A1(sum_ct[4]), .A2(n2868), .B1(n2869), .B2(ct[4]), .ZN(
        n2867) );
  INV_X1 U2159 ( .A(n2870), .ZN(n3357) );
  AOI22_X1 U2160 ( .A1(sum_ct[3]), .A2(n2868), .B1(n2869), .B2(ct[3]), .ZN(
        n2870) );
  INV_X1 U2161 ( .A(n2871), .ZN(n3358) );
  AOI22_X1 U2162 ( .A1(sum_ct[5]), .A2(n2868), .B1(n2869), .B2(ct[5]), .ZN(
        n2871) );
  INV_X1 U2163 ( .A(n2872), .ZN(n3359) );
  AOI22_X1 U2164 ( .A1(sum_ct[2]), .A2(n2868), .B1(n2869), .B2(ct[2]), .ZN(
        n2872) );
  INV_X1 U2165 ( .A(n2873), .ZN(n3360) );
  AOI22_X1 U2166 ( .A1(sum_ct[1]), .A2(n2868), .B1(n2869), .B2(ct[1]), .ZN(
        n2873) );
  INV_X1 U2167 ( .A(n2874), .ZN(n3361) );
  AOI22_X1 U2168 ( .A1(sum_ct[0]), .A2(n2868), .B1(n2869), .B2(ct[0]), .ZN(
        n2874) );
  AOI21_X1 U2169 ( .B1(n2875), .B2(n2876), .A(n2869), .ZN(n2868) );
  INV_X1 U2170 ( .A(n2877), .ZN(n2869) );
  OAI211_X1 U2171 ( .C1(n2878), .C2(n2876), .A(n2879), .B(n2875), .ZN(n2877)
         );
  OAI221_X1 U2172 ( .B1(n2880), .B2(n2836), .C1(n2881), .C2(n2882), .A(n2883), 
        .ZN(n999) );
  AOI22_X1 U2173 ( .A1(n2864), .A2(PR_1[11]), .B1(N275), .B2(n2884), .ZN(n2883) );
  INV_X1 U2174 ( .A(i_dividend[11]), .ZN(n2882) );
  OAI221_X1 U2175 ( .B1(n2880), .B2(n2837), .C1(n2881), .C2(n2885), .A(n2886), 
        .ZN(n998) );
  AOI22_X1 U2176 ( .A1(n2864), .A2(PR_1[12]), .B1(N276), .B2(n2884), .ZN(n2886) );
  INV_X1 U2177 ( .A(i_dividend[12]), .ZN(n2885) );
  OAI221_X1 U2178 ( .B1(n2880), .B2(n2838), .C1(n2881), .C2(n2887), .A(n2888), 
        .ZN(n997) );
  AOI22_X1 U2179 ( .A1(n2864), .A2(PR_1[13]), .B1(N277), .B2(n2884), .ZN(n2888) );
  INV_X1 U2180 ( .A(i_dividend[13]), .ZN(n2887) );
  OAI221_X1 U2181 ( .B1(n2880), .B2(n2839), .C1(n2881), .C2(n2889), .A(n2890), 
        .ZN(n996) );
  AOI22_X1 U2182 ( .A1(n2864), .A2(PR_1[14]), .B1(N278), .B2(n2884), .ZN(n2890) );
  INV_X1 U2183 ( .A(i_dividend[14]), .ZN(n2889) );
  OAI221_X1 U2184 ( .B1(n2880), .B2(n2840), .C1(n2881), .C2(n2891), .A(n2892), 
        .ZN(n995) );
  AOI22_X1 U2185 ( .A1(n2864), .A2(PR_1[15]), .B1(N279), .B2(n2884), .ZN(n2892) );
  INV_X1 U2186 ( .A(i_dividend[15]), .ZN(n2891) );
  OAI221_X1 U2187 ( .B1(n2880), .B2(n2841), .C1(n2881), .C2(n2893), .A(n2894), 
        .ZN(n994) );
  AOI22_X1 U2188 ( .A1(n2864), .A2(PR_1[16]), .B1(N280), .B2(n2884), .ZN(n2894) );
  INV_X1 U2189 ( .A(i_dividend[16]), .ZN(n2893) );
  OAI221_X1 U2190 ( .B1(n2880), .B2(n2842), .C1(n2881), .C2(n2895), .A(n2896), 
        .ZN(n993) );
  AOI22_X1 U2191 ( .A1(n2864), .A2(PR_1[17]), .B1(N281), .B2(n2884), .ZN(n2896) );
  INV_X1 U2192 ( .A(i_dividend[17]), .ZN(n2895) );
  OAI221_X1 U2193 ( .B1(n2880), .B2(n2843), .C1(n2881), .C2(n2897), .A(n2898), 
        .ZN(n992) );
  AOI22_X1 U2194 ( .A1(n2864), .A2(PR_1[18]), .B1(N282), .B2(n2884), .ZN(n2898) );
  INV_X1 U2195 ( .A(i_dividend[18]), .ZN(n2897) );
  OAI221_X1 U2196 ( .B1(n2880), .B2(n2844), .C1(n2881), .C2(n2899), .A(n2900), 
        .ZN(n991) );
  AOI22_X1 U2197 ( .A1(n2864), .A2(PR_1[19]), .B1(N283), .B2(n2884), .ZN(n2900) );
  INV_X1 U2198 ( .A(i_dividend[19]), .ZN(n2899) );
  OAI221_X1 U2199 ( .B1(n2880), .B2(n2845), .C1(n2881), .C2(n2901), .A(n2902), 
        .ZN(n990) );
  AOI22_X1 U2200 ( .A1(n2864), .A2(PR_1[20]), .B1(N284), .B2(n2884), .ZN(n2902) );
  INV_X1 U2201 ( .A(i_dividend[20]), .ZN(n2901) );
  OAI221_X1 U2202 ( .B1(n2880), .B2(n2846), .C1(n2881), .C2(n2903), .A(n2904), 
        .ZN(n989) );
  AOI22_X1 U2203 ( .A1(n2864), .A2(PR_1[21]), .B1(N285), .B2(n2884), .ZN(n2904) );
  INV_X1 U2204 ( .A(i_dividend[21]), .ZN(n2903) );
  OAI221_X1 U2205 ( .B1(n2880), .B2(n2818), .C1(n2881), .C2(n2905), .A(n2906), 
        .ZN(n988) );
  AOI22_X1 U2206 ( .A1(n2864), .A2(PR_1[22]), .B1(N286), .B2(n2884), .ZN(n2906) );
  INV_X1 U2207 ( .A(i_dividend[22]), .ZN(n2905) );
  OAI221_X1 U2208 ( .B1(n2880), .B2(n2819), .C1(n2881), .C2(n2907), .A(n2908), 
        .ZN(n987) );
  AOI22_X1 U2209 ( .A1(n2864), .A2(PR_1[23]), .B1(N287), .B2(n2884), .ZN(n2908) );
  INV_X1 U2210 ( .A(i_dividend[23]), .ZN(n2907) );
  OAI221_X1 U2211 ( .B1(n2880), .B2(n2820), .C1(n2881), .C2(n2909), .A(n2910), 
        .ZN(n986) );
  AOI22_X1 U2212 ( .A1(n2864), .A2(PR_1[24]), .B1(N288), .B2(n2884), .ZN(n2910) );
  INV_X1 U2213 ( .A(i_dividend[24]), .ZN(n2909) );
  OAI221_X1 U2214 ( .B1(n2880), .B2(n2824), .C1(n2881), .C2(n2911), .A(n2912), 
        .ZN(n985) );
  AOI22_X1 U2215 ( .A1(n2864), .A2(PR_1[25]), .B1(N289), .B2(n2884), .ZN(n2912) );
  INV_X1 U2216 ( .A(i_dividend[25]), .ZN(n2911) );
  OAI221_X1 U2217 ( .B1(n2880), .B2(n2815), .C1(n2881), .C2(n2913), .A(n2914), 
        .ZN(n984) );
  AOI22_X1 U2218 ( .A1(n2864), .A2(PR_1[26]), .B1(N290), .B2(n2884), .ZN(n2914) );
  INV_X1 U2219 ( .A(i_dividend[26]), .ZN(n2913) );
  OAI221_X1 U2220 ( .B1(n2880), .B2(n2821), .C1(n2881), .C2(n2915), .A(n2916), 
        .ZN(n983) );
  AOI22_X1 U2221 ( .A1(n2864), .A2(PR_1[27]), .B1(N291), .B2(n2884), .ZN(n2916) );
  INV_X1 U2222 ( .A(i_dividend[27]), .ZN(n2915) );
  OAI221_X1 U2223 ( .B1(n2880), .B2(n2822), .C1(n2881), .C2(n2917), .A(n2918), 
        .ZN(n982) );
  AOI22_X1 U2224 ( .A1(n2864), .A2(PR_1[28]), .B1(N292), .B2(n2884), .ZN(n2918) );
  INV_X1 U2225 ( .A(i_dividend[28]), .ZN(n2917) );
  OAI221_X1 U2226 ( .B1(n2880), .B2(n2823), .C1(n2881), .C2(n2919), .A(n2920), 
        .ZN(n981) );
  AOI22_X1 U2227 ( .A1(n2864), .A2(PR_1[29]), .B1(N293), .B2(n2884), .ZN(n2920) );
  INV_X1 U2228 ( .A(i_dividend[29]), .ZN(n2919) );
  OAI221_X1 U2229 ( .B1(n2880), .B2(n2816), .C1(n2881), .C2(n2921), .A(n2922), 
        .ZN(n980) );
  AOI22_X1 U2230 ( .A1(n2864), .A2(PR_1[30]), .B1(N294), .B2(n2884), .ZN(n2922) );
  INV_X1 U2231 ( .A(i_dividend[30]), .ZN(n2921) );
  OAI221_X1 U2232 ( .B1(n2880), .B2(n2814), .C1(n2881), .C2(n2923), .A(n2924), 
        .ZN(n979) );
  AOI22_X1 U2233 ( .A1(n2864), .A2(PR_1[31]), .B1(N295), .B2(n2884), .ZN(n2924) );
  INV_X1 U2234 ( .A(i_dividend[31]), .ZN(n2923) );
  OAI222_X1 U2235 ( .A1(n3307), .A2(n2925), .B1(n870), .B2(n2926), .C1(n2927), 
        .C2(n829), .ZN(n978) );
  MUX2_X1 U2236 ( .A(n3285), .B(sdata_o[6]), .S(n2866), .Z(n862) );
  MUX2_X1 U2237 ( .A(n3284), .B(sdata_o[7]), .S(n2866), .Z(n861) );
  MUX2_X1 U2238 ( .A(n3283), .B(sdata_o[8]), .S(n2866), .Z(n860) );
  MUX2_X1 U2239 ( .A(n3282), .B(sdata_o[9]), .S(n2866), .Z(n859) );
  MUX2_X1 U2240 ( .A(n3289), .B(sdata_o[10]), .S(n2866), .Z(n858) );
  MUX2_X1 U2241 ( .A(n3288), .B(sdata_o[11]), .S(n2866), .Z(n857) );
  MUX2_X1 U2242 ( .A(n3287), .B(sdata_o[12]), .S(n2866), .Z(n856) );
  MUX2_X1 U2243 ( .A(n3286), .B(sdata_o[13]), .S(n2866), .Z(n855) );
  MUX2_X1 U2244 ( .A(n3293), .B(sdata_o[14]), .S(n2866), .Z(n854) );
  MUX2_X1 U2245 ( .A(n3292), .B(sdata_o[15]), .S(n2866), .Z(n853) );
  MUX2_X1 U2246 ( .A(n3291), .B(sdata_o[16]), .S(n2866), .Z(n852) );
  MUX2_X1 U2247 ( .A(n3290), .B(sdata_o[17]), .S(n2866), .Z(n851) );
  MUX2_X1 U2248 ( .A(n3297), .B(sdata_o[18]), .S(n2866), .Z(n850) );
  MUX2_X1 U2249 ( .A(n3296), .B(sdata_o[19]), .S(n2866), .Z(n849) );
  MUX2_X1 U2250 ( .A(n3295), .B(sdata_o[20]), .S(n2866), .Z(n848) );
  MUX2_X1 U2251 ( .A(n3294), .B(sdata_o[21]), .S(n2866), .Z(n847) );
  MUX2_X1 U2252 ( .A(n3276), .B(sdata_o[22]), .S(n2866), .Z(n846) );
  MUX2_X1 U2253 ( .A(n3275), .B(sdata_o[23]), .S(n2866), .Z(n845) );
  MUX2_X1 U2254 ( .A(n3274), .B(sdata_o[24]), .S(n2866), .Z(n844) );
  MUX2_X1 U2255 ( .A(n3273), .B(sdata_o[25]), .S(n2866), .Z(n843) );
  MUX2_X1 U2256 ( .A(n3280), .B(sdata_o[26]), .S(n2866), .Z(n842) );
  MUX2_X1 U2257 ( .A(n3279), .B(sdata_o[27]), .S(n2866), .Z(n841) );
  MUX2_X1 U2258 ( .A(n3278), .B(sdata_o[28]), .S(n2866), .Z(n840) );
  MUX2_X1 U2259 ( .A(n3277), .B(sdata_o[29]), .S(n2866), .Z(n839) );
  MUX2_X1 U2260 ( .A(n3281), .B(sdata_o[30]), .S(n2866), .Z(n838) );
  INV_X1 U2261 ( .A(n2928), .ZN(n2786) );
  MUX2_X1 U2262 ( .A(n3304), .B(n3343), .S(n2929), .Z(n2928) );
  INV_X1 U2263 ( .A(n2930), .ZN(n2785) );
  MUX2_X1 U2264 ( .A(n3303), .B(n3344), .S(n2929), .Z(n2930) );
  INV_X1 U2265 ( .A(n2931), .ZN(n2784) );
  MUX2_X1 U2266 ( .A(n3302), .B(n3345), .S(n2929), .Z(n2931) );
  INV_X1 U2267 ( .A(n2932), .ZN(n2783) );
  MUX2_X1 U2268 ( .A(n3301), .B(n3346), .S(n2929), .Z(n2932) );
  OAI22_X1 U2269 ( .A1(n3305), .A2(n2927), .B1(n2880), .B2(n2933), .ZN(n1864)
         );
  OAI221_X1 U2270 ( .B1(n2925), .B2(n2788), .C1(n2927), .C2(n701), .A(n2934), 
        .ZN(n1297) );
  AOI222_X1 U2271 ( .A1(n2935), .A2(PR_1[30]), .B1(qp1[30]), .B2(n2863), .C1(
        q[30]), .C2(n2862), .ZN(n2934) );
  OAI221_X1 U2272 ( .B1(n2936), .B2(n2937), .C1(n2814), .C2(n2938), .A(n2939), 
        .ZN(n1296) );
  AOI222_X1 U2273 ( .A1(n2940), .A2(i_dividend[31]), .B1(n2941), .B2(
        sdata_o[31]), .C1(sum[31]), .C2(n2942), .ZN(n2939) );
  INV_X1 U2274 ( .A(i_divisor[31]), .ZN(n2937) );
  OAI211_X1 U2275 ( .C1(n941), .C2(n2927), .A(n2943), .B(n2881), .ZN(n1293) );
  OAI211_X1 U2276 ( .C1(n949), .C2(n2933), .A(n2944), .B(n2945), .ZN(n1292) );
  AOI222_X1 U2277 ( .A1(reg_b[0]), .A2(n2946), .B1(n2935), .B2(PR_1[0]), .C1(
        n2947), .C2(n3348), .ZN(n2945) );
  AOI22_X1 U2278 ( .A1(qp1[0]), .A2(n2863), .B1(q[0]), .B2(n2862), .ZN(n2944)
         );
  OAI211_X1 U2279 ( .C1(n948), .C2(n2933), .A(n2948), .B(n2949), .ZN(n1291) );
  AOI222_X1 U2280 ( .A1(reg_b[1]), .A2(n2946), .B1(n2935), .B2(PR_1[1]), .C1(
        n2947), .C2(n3342), .ZN(n2949) );
  AOI22_X1 U2281 ( .A1(qp1[1]), .A2(n2863), .B1(q[1]), .B2(n2862), .ZN(n2948)
         );
  OAI211_X1 U2282 ( .C1(n947), .C2(n2933), .A(n2950), .B(n2951), .ZN(n1290) );
  AOI222_X1 U2283 ( .A1(reg_b[2]), .A2(n2946), .B1(n2935), .B2(PR_1[2]), .C1(
        n2947), .C2(n3340), .ZN(n2951) );
  AOI22_X1 U2284 ( .A1(qp1[2]), .A2(n2863), .B1(q[2]), .B2(n2862), .ZN(n2950)
         );
  OAI211_X1 U2285 ( .C1(n946), .C2(n2933), .A(n2952), .B(n2953), .ZN(n1289) );
  AOI222_X1 U2286 ( .A1(reg_b[3]), .A2(n2946), .B1(n2935), .B2(PR_1[3]), .C1(
        n2947), .C2(n3338), .ZN(n2953) );
  AOI22_X1 U2287 ( .A1(qp1[3]), .A2(n2863), .B1(q[3]), .B2(n2862), .ZN(n2952)
         );
  OAI211_X1 U2288 ( .C1(n945), .C2(n2933), .A(n2954), .B(n2955), .ZN(n1288) );
  AOI222_X1 U2289 ( .A1(reg_b[4]), .A2(n2946), .B1(n2935), .B2(PR_1[4]), .C1(
        n2947), .C2(n3336), .ZN(n2955) );
  AOI22_X1 U2290 ( .A1(qp1[4]), .A2(n2863), .B1(q[4]), .B2(n2862), .ZN(n2954)
         );
  OAI211_X1 U2291 ( .C1(n944), .C2(n2933), .A(n2956), .B(n2957), .ZN(n1287) );
  AOI222_X1 U2292 ( .A1(reg_b[5]), .A2(n2946), .B1(n2935), .B2(PR_1[5]), .C1(
        n2947), .C2(n3334), .ZN(n2957) );
  AOI22_X1 U2293 ( .A1(qp1[5]), .A2(n2863), .B1(q[5]), .B2(n2862), .ZN(n2956)
         );
  OAI221_X1 U2294 ( .B1(n2925), .B2(n2787), .C1(n2927), .C2(n708), .A(n2958), 
        .ZN(n1286) );
  AOI222_X1 U2295 ( .A1(n2935), .A2(PR_1[6]), .B1(qp1[6]), .B2(n2863), .C1(
        q[6]), .C2(n2862), .ZN(n2958) );
  OAI221_X1 U2296 ( .B1(n2925), .B2(n2848), .C1(n2927), .C2(n709), .A(n2959), 
        .ZN(n1285) );
  AOI222_X1 U2297 ( .A1(n2935), .A2(PR_1[7]), .B1(qp1[7]), .B2(n2863), .C1(
        q[7]), .C2(n2862), .ZN(n2959) );
  OAI221_X1 U2298 ( .B1(n2925), .B2(n2801), .C1(n2927), .C2(n710), .A(n2960), 
        .ZN(n1284) );
  AOI222_X1 U2299 ( .A1(n2935), .A2(PR_1[8]), .B1(qp1[8]), .B2(n2863), .C1(
        q[8]), .C2(n2862), .ZN(n2960) );
  OAI221_X1 U2300 ( .B1(n2925), .B2(n2794), .C1(n2927), .C2(n711), .A(n2961), 
        .ZN(n1283) );
  AOI222_X1 U2301 ( .A1(n2935), .A2(PR_1[9]), .B1(qp1[9]), .B2(n2863), .C1(
        q[9]), .C2(n2862), .ZN(n2961) );
  OAI221_X1 U2302 ( .B1(n2925), .B2(n2792), .C1(n2927), .C2(n712), .A(n2962), 
        .ZN(n1282) );
  AOI222_X1 U2303 ( .A1(n2935), .A2(PR_1[10]), .B1(qp1[10]), .B2(n2863), .C1(
        q[10]), .C2(n2862), .ZN(n2962) );
  OAI221_X1 U2304 ( .B1(n2925), .B2(n2847), .C1(n2927), .C2(n713), .A(n2963), 
        .ZN(n1281) );
  AOI222_X1 U2305 ( .A1(n2935), .A2(PR_1[11]), .B1(qp1[11]), .B2(n2863), .C1(
        q[11]), .C2(n2862), .ZN(n2963) );
  OAI221_X1 U2306 ( .B1(n2925), .B2(n2800), .C1(n2927), .C2(n714), .A(n2964), 
        .ZN(n1280) );
  AOI222_X1 U2307 ( .A1(n2935), .A2(PR_1[12]), .B1(qp1[12]), .B2(n2863), .C1(
        q[12]), .C2(n2862), .ZN(n2964) );
  OAI221_X1 U2308 ( .B1(n2925), .B2(n2793), .C1(n2927), .C2(n715), .A(n2965), 
        .ZN(n1279) );
  AOI222_X1 U2309 ( .A1(n2935), .A2(PR_1[13]), .B1(qp1[13]), .B2(n2863), .C1(
        q[13]), .C2(n2862), .ZN(n2965) );
  OAI221_X1 U2310 ( .B1(n2925), .B2(n2791), .C1(n2927), .C2(n716), .A(n2966), 
        .ZN(n1278) );
  AOI222_X1 U2311 ( .A1(n2935), .A2(PR_1[14]), .B1(qp1[14]), .B2(n2863), .C1(
        q[14]), .C2(n2862), .ZN(n2966) );
  OAI221_X1 U2312 ( .B1(n2925), .B2(n2852), .C1(n2927), .C2(n717), .A(n2967), 
        .ZN(n1277) );
  AOI222_X1 U2313 ( .A1(n2935), .A2(PR_1[15]), .B1(qp1[15]), .B2(n2863), .C1(
        q[15]), .C2(n2862), .ZN(n2967) );
  OAI221_X1 U2314 ( .B1(n2925), .B2(n2805), .C1(n2927), .C2(n718), .A(n2968), 
        .ZN(n1276) );
  AOI222_X1 U2315 ( .A1(n2935), .A2(PR_1[16]), .B1(qp1[16]), .B2(n2863), .C1(
        q[16]), .C2(n2862), .ZN(n2968) );
  OAI221_X1 U2316 ( .B1(n2925), .B2(n2798), .C1(n2927), .C2(n719), .A(n2969), 
        .ZN(n1275) );
  AOI222_X1 U2317 ( .A1(n2935), .A2(PR_1[17]), .B1(qp1[17]), .B2(n2863), .C1(
        q[17]), .C2(n2862), .ZN(n2969) );
  OAI221_X1 U2318 ( .B1(n2925), .B2(n2858), .C1(n2927), .C2(n720), .A(n2970), 
        .ZN(n1274) );
  AOI222_X1 U2319 ( .A1(n2935), .A2(PR_1[18]), .B1(qp1[18]), .B2(n2863), .C1(
        q[18]), .C2(n2862), .ZN(n2970) );
  OAI221_X1 U2320 ( .B1(n2925), .B2(n2851), .C1(n2927), .C2(n721), .A(n2971), 
        .ZN(n1273) );
  AOI222_X1 U2321 ( .A1(n2935), .A2(PR_1[19]), .B1(qp1[19]), .B2(n2863), .C1(
        q[19]), .C2(n2862), .ZN(n2971) );
  OAI221_X1 U2322 ( .B1(n2925), .B2(n2804), .C1(n2927), .C2(n722), .A(n2972), 
        .ZN(n1272) );
  AOI222_X1 U2323 ( .A1(n2935), .A2(PR_1[20]), .B1(qp1[20]), .B2(n2863), .C1(
        q[20]), .C2(n2862), .ZN(n2972) );
  OAI221_X1 U2324 ( .B1(n2925), .B2(n2797), .C1(n2927), .C2(n723), .A(n2973), 
        .ZN(n1271) );
  AOI222_X1 U2325 ( .A1(n2935), .A2(PR_1[21]), .B1(qp1[21]), .B2(n2863), .C1(
        q[21]), .C2(n2862), .ZN(n2973) );
  OAI221_X1 U2326 ( .B1(n2925), .B2(n2850), .C1(n2927), .C2(n724), .A(n2974), 
        .ZN(n1270) );
  AOI222_X1 U2327 ( .A1(n2935), .A2(PR_1[22]), .B1(qp1[22]), .B2(n2863), .C1(
        q[22]), .C2(n2862), .ZN(n2974) );
  OAI221_X1 U2328 ( .B1(n2925), .B2(n2803), .C1(n2927), .C2(n725), .A(n2975), 
        .ZN(n1269) );
  AOI222_X1 U2329 ( .A1(n2935), .A2(PR_1[23]), .B1(qp1[23]), .B2(n2863), .C1(
        q[23]), .C2(n2862), .ZN(n2975) );
  OAI221_X1 U2330 ( .B1(n2925), .B2(n2796), .C1(n2927), .C2(n726), .A(n2976), 
        .ZN(n1268) );
  AOI222_X1 U2331 ( .A1(n2935), .A2(PR_1[24]), .B1(qp1[24]), .B2(n2863), .C1(
        q[24]), .C2(n2862), .ZN(n2976) );
  OAI221_X1 U2332 ( .B1(n2925), .B2(n2790), .C1(n2927), .C2(n727), .A(n2977), 
        .ZN(n1267) );
  AOI222_X1 U2333 ( .A1(n2935), .A2(PR_1[25]), .B1(qp1[25]), .B2(n2863), .C1(
        q[25]), .C2(n2862), .ZN(n2977) );
  OAI221_X1 U2334 ( .B1(n2925), .B2(n2849), .C1(n2927), .C2(n728), .A(n2978), 
        .ZN(n1266) );
  AOI222_X1 U2335 ( .A1(n2935), .A2(PR_1[26]), .B1(qp1[26]), .B2(n2863), .C1(
        q[26]), .C2(n2862), .ZN(n2978) );
  OAI221_X1 U2336 ( .B1(n2925), .B2(n2802), .C1(n2927), .C2(n729), .A(n2979), 
        .ZN(n1265) );
  AOI222_X1 U2337 ( .A1(n2935), .A2(PR_1[27]), .B1(qp1[27]), .B2(n2863), .C1(
        q[27]), .C2(n2862), .ZN(n2979) );
  OAI221_X1 U2338 ( .B1(n2925), .B2(n2795), .C1(n2927), .C2(n730), .A(n2980), 
        .ZN(n1264) );
  AOI222_X1 U2339 ( .A1(n2935), .A2(PR_1[28]), .B1(qp1[28]), .B2(n2863), .C1(
        q[28]), .C2(n2862), .ZN(n2980) );
  OAI221_X1 U2340 ( .B1(n2925), .B2(n2789), .C1(n2927), .C2(n731), .A(n2981), 
        .ZN(n1263) );
  AOI222_X1 U2341 ( .A1(n2935), .A2(PR_1[29]), .B1(qp1[29]), .B2(n2863), .C1(
        q[29]), .C2(n2862), .ZN(n2981) );
  MUX2_X1 U2342 ( .A(sum[0]), .B(o_remainder[0]), .S(n2985), .Z(n1262) );
  MUX2_X1 U2343 ( .A(sum[1]), .B(o_remainder[1]), .S(n2985), .Z(n1261) );
  MUX2_X1 U2344 ( .A(sum[2]), .B(o_remainder[2]), .S(n2985), .Z(n1260) );
  MUX2_X1 U2345 ( .A(sum[3]), .B(o_remainder[3]), .S(n2985), .Z(n1259) );
  MUX2_X1 U2346 ( .A(sum[4]), .B(o_remainder[4]), .S(n2985), .Z(n1258) );
  MUX2_X1 U2347 ( .A(sum[5]), .B(o_remainder[5]), .S(n2985), .Z(n1257) );
  MUX2_X1 U2348 ( .A(sum[6]), .B(o_remainder[6]), .S(n2985), .Z(n1256) );
  MUX2_X1 U2349 ( .A(sum[7]), .B(o_remainder[7]), .S(n2985), .Z(n1255) );
  MUX2_X1 U2350 ( .A(sum[8]), .B(o_remainder[8]), .S(n2985), .Z(n1254) );
  MUX2_X1 U2351 ( .A(sum[9]), .B(o_remainder[9]), .S(n2985), .Z(n1253) );
  MUX2_X1 U2352 ( .A(sum[10]), .B(o_remainder[10]), .S(n2985), .Z(n1252) );
  MUX2_X1 U2353 ( .A(sum[11]), .B(o_remainder[11]), .S(n2985), .Z(n1251) );
  MUX2_X1 U2354 ( .A(sum[12]), .B(o_remainder[12]), .S(n2985), .Z(n1250) );
  MUX2_X1 U2355 ( .A(sum[13]), .B(o_remainder[13]), .S(n2985), .Z(n1249) );
  MUX2_X1 U2356 ( .A(sum[14]), .B(o_remainder[14]), .S(n2985), .Z(n1248) );
  MUX2_X1 U2357 ( .A(sum[15]), .B(o_remainder[15]), .S(n2985), .Z(n1247) );
  MUX2_X1 U2358 ( .A(sum[16]), .B(o_remainder[16]), .S(n2985), .Z(n1246) );
  MUX2_X1 U2359 ( .A(sum[17]), .B(o_remainder[17]), .S(n2985), .Z(n1245) );
  MUX2_X1 U2360 ( .A(sum[18]), .B(o_remainder[18]), .S(n2985), .Z(n1244) );
  MUX2_X1 U2361 ( .A(sum[19]), .B(o_remainder[19]), .S(n2985), .Z(n1243) );
  MUX2_X1 U2362 ( .A(sum[20]), .B(o_remainder[20]), .S(n2985), .Z(n1242) );
  MUX2_X1 U2363 ( .A(sum[21]), .B(o_remainder[21]), .S(n2985), .Z(n1241) );
  MUX2_X1 U2364 ( .A(sum[22]), .B(o_remainder[22]), .S(n2985), .Z(n1240) );
  MUX2_X1 U2365 ( .A(sum[23]), .B(o_remainder[23]), .S(n2985), .Z(n1239) );
  MUX2_X1 U2366 ( .A(sum[24]), .B(o_remainder[24]), .S(n2985), .Z(n1238) );
  MUX2_X1 U2367 ( .A(sum[25]), .B(o_remainder[25]), .S(n2985), .Z(n1237) );
  MUX2_X1 U2368 ( .A(sum[26]), .B(o_remainder[26]), .S(n2985), .Z(n1236) );
  MUX2_X1 U2369 ( .A(sum[27]), .B(o_remainder[27]), .S(n2985), .Z(n1235) );
  MUX2_X1 U2370 ( .A(sum[28]), .B(o_remainder[28]), .S(n2985), .Z(n1234) );
  MUX2_X1 U2371 ( .A(sum[29]), .B(o_remainder[29]), .S(n2985), .Z(n1233) );
  MUX2_X1 U2372 ( .A(sum[30]), .B(o_remainder[30]), .S(n2985), .Z(n1232) );
  MUX2_X1 U2373 ( .A(sum[31]), .B(o_remainder[31]), .S(n2985), .Z(n1231) );
  NAND2_X1 U2374 ( .A1(n2865), .A2(n2985), .ZN(n1230) );
  NAND2_X1 U2375 ( .A1(ready), .A2(i_start), .ZN(n2865) );
  MUX2_X1 U2376 ( .A(n2986), .B(state[5]), .S(n2987), .Z(n1229) );
  MUX2_X1 U2377 ( .A(n2988), .B(state[1]), .S(n2987), .Z(n1228) );
  MUX2_X1 U2378 ( .A(n3272), .B(i_dividend[31]), .S(n2989), .Z(n1227) );
  MUX2_X1 U2379 ( .A(n2990), .B(state[2]), .S(n2987), .Z(n1226) );
  MUX2_X1 U2380 ( .A(n2991), .B(state[3]), .S(n2987), .Z(n1225) );
  MUX2_X1 U2381 ( .A(o_quotient[0]), .B(sum[0]), .S(n2884), .Z(n1224) );
  MUX2_X1 U2382 ( .A(o_quotient[1]), .B(sum[1]), .S(n2884), .Z(n1223) );
  MUX2_X1 U2383 ( .A(o_quotient[2]), .B(sum[2]), .S(n2884), .Z(n1222) );
  MUX2_X1 U2384 ( .A(o_quotient[3]), .B(sum[3]), .S(n2884), .Z(n1221) );
  MUX2_X1 U2385 ( .A(o_quotient[4]), .B(sum[4]), .S(n2884), .Z(n1220) );
  MUX2_X1 U2386 ( .A(o_quotient[5]), .B(sum[5]), .S(n2884), .Z(n1219) );
  MUX2_X1 U2387 ( .A(o_quotient[6]), .B(sum[6]), .S(n2884), .Z(n1218) );
  MUX2_X1 U2388 ( .A(o_quotient[7]), .B(sum[7]), .S(n2884), .Z(n1217) );
  MUX2_X1 U2389 ( .A(o_quotient[8]), .B(sum[8]), .S(n2884), .Z(n1216) );
  MUX2_X1 U2390 ( .A(o_quotient[9]), .B(sum[9]), .S(n2884), .Z(n1215) );
  MUX2_X1 U2391 ( .A(o_quotient[10]), .B(sum[10]), .S(n2884), .Z(n1214) );
  MUX2_X1 U2392 ( .A(o_quotient[11]), .B(sum[11]), .S(n2884), .Z(n1213) );
  MUX2_X1 U2393 ( .A(o_quotient[12]), .B(sum[12]), .S(n2884), .Z(n1212) );
  MUX2_X1 U2394 ( .A(o_quotient[13]), .B(sum[13]), .S(n2884), .Z(n1211) );
  MUX2_X1 U2395 ( .A(o_quotient[14]), .B(sum[14]), .S(n2884), .Z(n1210) );
  MUX2_X1 U2396 ( .A(o_quotient[15]), .B(sum[15]), .S(n2884), .Z(n1209) );
  MUX2_X1 U2397 ( .A(o_quotient[16]), .B(sum[16]), .S(n2884), .Z(n1208) );
  MUX2_X1 U2398 ( .A(o_quotient[17]), .B(sum[17]), .S(n2884), .Z(n1207) );
  MUX2_X1 U2399 ( .A(o_quotient[18]), .B(sum[18]), .S(n2884), .Z(n1206) );
  MUX2_X1 U2400 ( .A(o_quotient[19]), .B(sum[19]), .S(n2884), .Z(n1205) );
  MUX2_X1 U2401 ( .A(o_quotient[20]), .B(sum[20]), .S(n2884), .Z(n1204) );
  MUX2_X1 U2402 ( .A(o_quotient[21]), .B(sum[21]), .S(n2884), .Z(n1203) );
  MUX2_X1 U2403 ( .A(o_quotient[22]), .B(sum[22]), .S(n2884), .Z(n1202) );
  MUX2_X1 U2404 ( .A(o_quotient[23]), .B(sum[23]), .S(n2884), .Z(n1201) );
  MUX2_X1 U2405 ( .A(o_quotient[24]), .B(sum[24]), .S(n2884), .Z(n1200) );
  MUX2_X1 U2406 ( .A(o_quotient[25]), .B(sum[25]), .S(n2884), .Z(n1199) );
  MUX2_X1 U2407 ( .A(o_quotient[26]), .B(sum[26]), .S(n2884), .Z(n1198) );
  MUX2_X1 U2408 ( .A(o_quotient[27]), .B(sum[27]), .S(n2884), .Z(n1197) );
  MUX2_X1 U2409 ( .A(o_quotient[28]), .B(sum[28]), .S(n2884), .Z(n1196) );
  MUX2_X1 U2410 ( .A(o_quotient[29]), .B(sum[29]), .S(n2884), .Z(n1195) );
  MUX2_X1 U2411 ( .A(o_quotient[30]), .B(sum[30]), .S(n2884), .Z(n1194) );
  MUX2_X1 U2412 ( .A(o_quotient[31]), .B(sum[31]), .S(n2884), .Z(n1193) );
  MUX2_X1 U2413 ( .A(n2992), .B(state[4]), .S(n2987), .Z(n1192) );
  MUX2_X1 U2414 ( .A(n2993), .B(state[0]), .S(n2987), .Z(n1191) );
  AND4_X1 U2415 ( .A1(n2994), .A2(n2995), .A3(n2996), .A4(n2985), .ZN(n2987)
         );
  NOR2_X1 U2416 ( .A1(n977), .A2(n2989), .ZN(n2996) );
  NAND2_X1 U2417 ( .A1(n2997), .A2(n2879), .ZN(n977) );
  NAND3_X1 U2418 ( .A1(n2998), .A2(ct[5]), .A3(n2991), .ZN(n2879) );
  OAI21_X1 U2419 ( .B1(n3346), .B2(n2999), .A(n3000), .ZN(n1190) );
  NAND2_X1 U2420 ( .A1(shifted_o[0]), .A2(n3001), .ZN(n3000) );
  OAI21_X1 U2421 ( .B1(n3345), .B2(n2999), .A(n3002), .ZN(n1189) );
  NAND2_X1 U2422 ( .A1(shifted_o[1]), .A2(n3001), .ZN(n3002) );
  OAI21_X1 U2423 ( .B1(n3344), .B2(n2999), .A(n3003), .ZN(n1188) );
  NAND2_X1 U2424 ( .A1(shifted_o[2]), .A2(n3001), .ZN(n3003) );
  OAI21_X1 U2425 ( .B1(n3343), .B2(n2999), .A(n3004), .ZN(n1187) );
  NAND2_X1 U2426 ( .A1(shifted_o[3]), .A2(n3001), .ZN(n3004) );
  NAND2_X1 U2427 ( .A1(n3005), .A2(n2995), .ZN(n2999) );
  INV_X1 U2428 ( .A(n3001), .ZN(n3005) );
  NAND2_X1 U2429 ( .A1(n2875), .A2(n2880), .ZN(n3001) );
  OAI221_X1 U2430 ( .B1(n2936), .B2(n3006), .C1(n2938), .C2(n2825), .A(n3007), 
        .ZN(n1186) );
  AOI222_X1 U2431 ( .A1(i_dividend[0]), .A2(n2940), .B1(n2941), .B2(sdata_o[0]), .C1(sum[0]), .C2(n2942), .ZN(n3007) );
  INV_X1 U2432 ( .A(i_divisor[0]), .ZN(n3006) );
  OAI221_X1 U2433 ( .B1(n2936), .B2(n3008), .C1(n2938), .C2(n2826), .A(n3009), 
        .ZN(n1185) );
  AOI222_X1 U2434 ( .A1(i_dividend[1]), .A2(n2940), .B1(n2941), .B2(sdata_o[1]), .C1(sum[1]), .C2(n2942), .ZN(n3009) );
  INV_X1 U2435 ( .A(i_divisor[1]), .ZN(n3008) );
  OAI221_X1 U2436 ( .B1(n2936), .B2(n3010), .C1(n2938), .C2(n2827), .A(n3011), 
        .ZN(n1184) );
  AOI222_X1 U2437 ( .A1(i_dividend[2]), .A2(n2940), .B1(n2941), .B2(sdata_o[2]), .C1(sum[2]), .C2(n2942), .ZN(n3011) );
  INV_X1 U2438 ( .A(i_divisor[2]), .ZN(n3010) );
  OAI221_X1 U2439 ( .B1(n2936), .B2(n3012), .C1(n2938), .C2(n2828), .A(n3013), 
        .ZN(n1183) );
  AOI222_X1 U2440 ( .A1(i_dividend[3]), .A2(n2940), .B1(n2941), .B2(sdata_o[3]), .C1(sum[3]), .C2(n2942), .ZN(n3013) );
  INV_X1 U2441 ( .A(i_divisor[3]), .ZN(n3012) );
  OAI221_X1 U2442 ( .B1(n2936), .B2(n3014), .C1(n2938), .C2(n2829), .A(n3015), 
        .ZN(n1182) );
  AOI222_X1 U2443 ( .A1(i_dividend[4]), .A2(n2940), .B1(n2941), .B2(sdata_o[4]), .C1(sum[4]), .C2(n2942), .ZN(n3015) );
  INV_X1 U2444 ( .A(i_divisor[4]), .ZN(n3014) );
  OAI221_X1 U2445 ( .B1(n2936), .B2(n3016), .C1(n2938), .C2(n2830), .A(n3017), 
        .ZN(n1181) );
  AOI222_X1 U2446 ( .A1(i_dividend[5]), .A2(n2940), .B1(n2941), .B2(sdata_o[5]), .C1(sum[5]), .C2(n2942), .ZN(n3017) );
  INV_X1 U2447 ( .A(i_divisor[5]), .ZN(n3016) );
  OAI221_X1 U2448 ( .B1(n2936), .B2(n3018), .C1(n2938), .C2(n2831), .A(n3019), 
        .ZN(n1180) );
  AOI222_X1 U2449 ( .A1(i_dividend[6]), .A2(n2940), .B1(n2941), .B2(sdata_o[6]), .C1(sum[6]), .C2(n2942), .ZN(n3019) );
  INV_X1 U2450 ( .A(i_divisor[6]), .ZN(n3018) );
  OAI221_X1 U2451 ( .B1(n2936), .B2(n3020), .C1(n2938), .C2(n2832), .A(n3021), 
        .ZN(n1179) );
  AOI222_X1 U2452 ( .A1(i_dividend[7]), .A2(n2940), .B1(n2941), .B2(sdata_o[7]), .C1(sum[7]), .C2(n2942), .ZN(n3021) );
  INV_X1 U2453 ( .A(i_divisor[7]), .ZN(n3020) );
  OAI221_X1 U2454 ( .B1(n2936), .B2(n3022), .C1(n2938), .C2(n2833), .A(n3023), 
        .ZN(n1178) );
  AOI222_X1 U2455 ( .A1(i_dividend[8]), .A2(n2940), .B1(n2941), .B2(sdata_o[8]), .C1(sum[8]), .C2(n2942), .ZN(n3023) );
  INV_X1 U2456 ( .A(i_divisor[8]), .ZN(n3022) );
  OAI221_X1 U2457 ( .B1(n2936), .B2(n3024), .C1(n2938), .C2(n2834), .A(n3025), 
        .ZN(n1177) );
  AOI222_X1 U2458 ( .A1(i_dividend[9]), .A2(n2940), .B1(n2941), .B2(sdata_o[9]), .C1(sum[9]), .C2(n2942), .ZN(n3025) );
  INV_X1 U2459 ( .A(i_divisor[9]), .ZN(n3024) );
  OAI221_X1 U2460 ( .B1(n2936), .B2(n3026), .C1(n2938), .C2(n2835), .A(n3027), 
        .ZN(n1176) );
  AOI222_X1 U2461 ( .A1(i_dividend[10]), .A2(n2940), .B1(n2941), .B2(
        sdata_o[10]), .C1(sum[10]), .C2(n2942), .ZN(n3027) );
  INV_X1 U2462 ( .A(i_divisor[10]), .ZN(n3026) );
  OAI221_X1 U2463 ( .B1(n2936), .B2(n3028), .C1(n2836), .C2(n2938), .A(n3029), 
        .ZN(n1175) );
  AOI222_X1 U2464 ( .A1(n2940), .A2(i_dividend[11]), .B1(n2941), .B2(
        sdata_o[11]), .C1(sum[11]), .C2(n2942), .ZN(n3029) );
  INV_X1 U2465 ( .A(i_divisor[11]), .ZN(n3028) );
  OAI221_X1 U2466 ( .B1(n2936), .B2(n3030), .C1(n2837), .C2(n2938), .A(n3031), 
        .ZN(n1174) );
  AOI222_X1 U2467 ( .A1(n2940), .A2(i_dividend[12]), .B1(n2941), .B2(
        sdata_o[12]), .C1(sum[12]), .C2(n2942), .ZN(n3031) );
  INV_X1 U2468 ( .A(i_divisor[12]), .ZN(n3030) );
  OAI221_X1 U2469 ( .B1(n2936), .B2(n3032), .C1(n2838), .C2(n2938), .A(n3033), 
        .ZN(n1173) );
  AOI222_X1 U2470 ( .A1(n2940), .A2(i_dividend[13]), .B1(n2941), .B2(
        sdata_o[13]), .C1(sum[13]), .C2(n2942), .ZN(n3033) );
  INV_X1 U2471 ( .A(i_divisor[13]), .ZN(n3032) );
  OAI221_X1 U2472 ( .B1(n2936), .B2(n3034), .C1(n2839), .C2(n2938), .A(n3035), 
        .ZN(n1172) );
  AOI222_X1 U2473 ( .A1(n2940), .A2(i_dividend[14]), .B1(n2941), .B2(
        sdata_o[14]), .C1(sum[14]), .C2(n2942), .ZN(n3035) );
  INV_X1 U2474 ( .A(i_divisor[14]), .ZN(n3034) );
  OAI221_X1 U2475 ( .B1(n2936), .B2(n3036), .C1(n2840), .C2(n2938), .A(n3037), 
        .ZN(n1171) );
  AOI222_X1 U2476 ( .A1(n2940), .A2(i_dividend[15]), .B1(n2941), .B2(
        sdata_o[15]), .C1(sum[15]), .C2(n2942), .ZN(n3037) );
  INV_X1 U2477 ( .A(i_divisor[15]), .ZN(n3036) );
  OAI221_X1 U2478 ( .B1(n2936), .B2(n3038), .C1(n2841), .C2(n2938), .A(n3039), 
        .ZN(n1170) );
  AOI222_X1 U2479 ( .A1(n2940), .A2(i_dividend[16]), .B1(n2941), .B2(
        sdata_o[16]), .C1(sum[16]), .C2(n2942), .ZN(n3039) );
  INV_X1 U2480 ( .A(i_divisor[16]), .ZN(n3038) );
  OAI221_X1 U2481 ( .B1(n2936), .B2(n3040), .C1(n2842), .C2(n2938), .A(n3041), 
        .ZN(n1169) );
  AOI222_X1 U2482 ( .A1(n2940), .A2(i_dividend[17]), .B1(n2941), .B2(
        sdata_o[17]), .C1(sum[17]), .C2(n2942), .ZN(n3041) );
  INV_X1 U2483 ( .A(i_divisor[17]), .ZN(n3040) );
  OAI221_X1 U2484 ( .B1(n2936), .B2(n3042), .C1(n2843), .C2(n2938), .A(n3043), 
        .ZN(n1168) );
  AOI222_X1 U2485 ( .A1(n2940), .A2(i_dividend[18]), .B1(n2941), .B2(
        sdata_o[18]), .C1(sum[18]), .C2(n2942), .ZN(n3043) );
  INV_X1 U2486 ( .A(i_divisor[18]), .ZN(n3042) );
  OAI221_X1 U2487 ( .B1(n2936), .B2(n3044), .C1(n2844), .C2(n2938), .A(n3045), 
        .ZN(n1167) );
  AOI222_X1 U2488 ( .A1(n2940), .A2(i_dividend[19]), .B1(n2941), .B2(
        sdata_o[19]), .C1(sum[19]), .C2(n2942), .ZN(n3045) );
  INV_X1 U2489 ( .A(i_divisor[19]), .ZN(n3044) );
  OAI221_X1 U2490 ( .B1(n2936), .B2(n3046), .C1(n2845), .C2(n2938), .A(n3047), 
        .ZN(n1166) );
  AOI222_X1 U2491 ( .A1(n2940), .A2(i_dividend[20]), .B1(n2941), .B2(
        sdata_o[20]), .C1(sum[20]), .C2(n2942), .ZN(n3047) );
  INV_X1 U2492 ( .A(i_divisor[20]), .ZN(n3046) );
  OAI221_X1 U2493 ( .B1(n2936), .B2(n3048), .C1(n2846), .C2(n2938), .A(n3049), 
        .ZN(n1165) );
  AOI222_X1 U2494 ( .A1(n2940), .A2(i_dividend[21]), .B1(n2941), .B2(
        sdata_o[21]), .C1(sum[21]), .C2(n2942), .ZN(n3049) );
  INV_X1 U2495 ( .A(i_divisor[21]), .ZN(n3048) );
  OAI221_X1 U2496 ( .B1(n2936), .B2(n3050), .C1(n2818), .C2(n2938), .A(n3051), 
        .ZN(n1164) );
  AOI222_X1 U2497 ( .A1(n2940), .A2(i_dividend[22]), .B1(n2941), .B2(
        sdata_o[22]), .C1(sum[22]), .C2(n2942), .ZN(n3051) );
  INV_X1 U2498 ( .A(i_divisor[22]), .ZN(n3050) );
  OAI221_X1 U2499 ( .B1(n2936), .B2(n3052), .C1(n2819), .C2(n2938), .A(n3053), 
        .ZN(n1163) );
  AOI222_X1 U2500 ( .A1(n2940), .A2(i_dividend[23]), .B1(n2941), .B2(
        sdata_o[23]), .C1(sum[23]), .C2(n2942), .ZN(n3053) );
  INV_X1 U2501 ( .A(i_divisor[23]), .ZN(n3052) );
  OAI221_X1 U2502 ( .B1(n2936), .B2(n3054), .C1(n2820), .C2(n2938), .A(n3055), 
        .ZN(n1162) );
  AOI222_X1 U2503 ( .A1(n2940), .A2(i_dividend[24]), .B1(n2941), .B2(
        sdata_o[24]), .C1(sum[24]), .C2(n2942), .ZN(n3055) );
  INV_X1 U2504 ( .A(i_divisor[24]), .ZN(n3054) );
  OAI221_X1 U2505 ( .B1(n2936), .B2(n3056), .C1(n2824), .C2(n2938), .A(n3057), 
        .ZN(n1161) );
  AOI222_X1 U2506 ( .A1(n2940), .A2(i_dividend[25]), .B1(n2941), .B2(
        sdata_o[25]), .C1(sum[25]), .C2(n2942), .ZN(n3057) );
  INV_X1 U2507 ( .A(i_divisor[25]), .ZN(n3056) );
  OAI221_X1 U2508 ( .B1(n2936), .B2(n3058), .C1(n2815), .C2(n2938), .A(n3059), 
        .ZN(n1160) );
  AOI222_X1 U2509 ( .A1(n2940), .A2(i_dividend[26]), .B1(n2941), .B2(
        sdata_o[26]), .C1(sum[26]), .C2(n2942), .ZN(n3059) );
  INV_X1 U2510 ( .A(i_divisor[26]), .ZN(n3058) );
  OAI221_X1 U2511 ( .B1(n2936), .B2(n3060), .C1(n2821), .C2(n2938), .A(n3061), 
        .ZN(n1159) );
  AOI222_X1 U2512 ( .A1(n2940), .A2(i_dividend[27]), .B1(n2941), .B2(
        sdata_o[27]), .C1(sum[27]), .C2(n2942), .ZN(n3061) );
  INV_X1 U2513 ( .A(i_divisor[27]), .ZN(n3060) );
  OAI221_X1 U2514 ( .B1(n2936), .B2(n3062), .C1(n2822), .C2(n2938), .A(n3063), 
        .ZN(n1158) );
  AOI222_X1 U2515 ( .A1(n2940), .A2(i_dividend[28]), .B1(n2941), .B2(
        sdata_o[28]), .C1(sum[28]), .C2(n2942), .ZN(n3063) );
  INV_X1 U2516 ( .A(i_divisor[28]), .ZN(n3062) );
  OAI221_X1 U2517 ( .B1(n2936), .B2(n3064), .C1(n2823), .C2(n2938), .A(n3065), 
        .ZN(n1157) );
  AOI222_X1 U2518 ( .A1(n2940), .A2(i_dividend[29]), .B1(n2941), .B2(
        sdata_o[29]), .C1(sum[29]), .C2(n2942), .ZN(n3065) );
  INV_X1 U2519 ( .A(i_divisor[29]), .ZN(n3064) );
  OAI221_X1 U2520 ( .B1(n2936), .B2(n3066), .C1(n2816), .C2(n2938), .A(n3067), 
        .ZN(n1156) );
  AOI222_X1 U2521 ( .A1(n2940), .A2(i_dividend[30]), .B1(n2941), .B2(
        sdata_o[30]), .C1(sum[30]), .C2(n2942), .ZN(n3067) );
  INV_X1 U2522 ( .A(i_divisor[30]), .ZN(n3066) );
  MUX2_X1 U2523 ( .A(sdata[0]), .B(n3306), .S(n2994), .Z(n1155) );
  MUX2_X1 U2524 ( .A(sdata[1]), .B(n3341), .S(n2994), .Z(n1154) );
  MUX2_X1 U2525 ( .A(sdata[2]), .B(n3339), .S(n2994), .Z(n1153) );
  MUX2_X1 U2526 ( .A(sdata[3]), .B(n3337), .S(n2994), .Z(n1152) );
  MUX2_X1 U2527 ( .A(sdata[4]), .B(n3335), .S(n2994), .Z(n1151) );
  MUX2_X1 U2528 ( .A(sdata[5]), .B(n3333), .S(n2994), .Z(n1150) );
  MUX2_X1 U2529 ( .A(sdata[6]), .B(n3332), .S(n2994), .Z(n1149) );
  MUX2_X1 U2530 ( .A(sdata[7]), .B(n3331), .S(n2994), .Z(n1148) );
  MUX2_X1 U2531 ( .A(sdata[8]), .B(n3330), .S(n2994), .Z(n1147) );
  MUX2_X1 U2532 ( .A(sdata[9]), .B(n3329), .S(n2994), .Z(n1146) );
  MUX2_X1 U2533 ( .A(sdata[10]), .B(n3328), .S(n2994), .Z(n1145) );
  MUX2_X1 U2534 ( .A(sdata[11]), .B(n3327), .S(n2994), .Z(n1144) );
  MUX2_X1 U2535 ( .A(sdata[12]), .B(n3326), .S(n2994), .Z(n1143) );
  MUX2_X1 U2536 ( .A(sdata[13]), .B(n3325), .S(n2994), .Z(n1142) );
  MUX2_X1 U2537 ( .A(sdata[14]), .B(n3324), .S(n2994), .Z(n1141) );
  MUX2_X1 U2538 ( .A(sdata[15]), .B(n3323), .S(n2994), .Z(n1140) );
  MUX2_X1 U2539 ( .A(sdata[16]), .B(n3322), .S(n2994), .Z(n1139) );
  MUX2_X1 U2540 ( .A(sdata[17]), .B(n3321), .S(n2994), .Z(n1138) );
  MUX2_X1 U2541 ( .A(sdata[18]), .B(n3320), .S(n2994), .Z(n1137) );
  MUX2_X1 U2542 ( .A(sdata[19]), .B(n3319), .S(n2994), .Z(n1136) );
  MUX2_X1 U2543 ( .A(sdata[20]), .B(n3318), .S(n2994), .Z(n1135) );
  MUX2_X1 U2544 ( .A(sdata[21]), .B(n3317), .S(n2994), .Z(n1134) );
  MUX2_X1 U2545 ( .A(sdata[22]), .B(n3316), .S(n2994), .Z(n1133) );
  MUX2_X1 U2546 ( .A(sdata[23]), .B(n3315), .S(n2994), .Z(n1132) );
  MUX2_X1 U2547 ( .A(sdata[24]), .B(n3314), .S(n2994), .Z(n1131) );
  MUX2_X1 U2548 ( .A(sdata[25]), .B(n3313), .S(n2994), .Z(n1130) );
  MUX2_X1 U2549 ( .A(sdata[26]), .B(n3312), .S(n2994), .Z(n1129) );
  MUX2_X1 U2550 ( .A(sdata[27]), .B(n3311), .S(n2994), .Z(n1128) );
  MUX2_X1 U2551 ( .A(sdata[28]), .B(n3310), .S(n2994), .Z(n1127) );
  MUX2_X1 U2552 ( .A(sdata[29]), .B(n3309), .S(n2994), .Z(n1126) );
  MUX2_X1 U2553 ( .A(sdata[30]), .B(n3308), .S(n2994), .Z(n1125) );
  MUX2_X1 U2554 ( .A(sdata[31]), .B(n3299), .S(n2994), .Z(n1124) );
  XOR2_X1 U2555 ( .A(n2814), .B(sdata[30]), .Z(n3068) );
  NAND2_X1 U2556 ( .A1(n2998), .A2(n2988), .ZN(n2875) );
  AND4_X1 U2557 ( .A1(n3069), .A2(state[5]), .A3(n2853), .A4(n2806), .ZN(n2988) );
  MUX2_X1 U2558 ( .A(n2998), .B(n3298), .S(n3070), .Z(n1113) );
  NOR2_X1 U2559 ( .A1(n2929), .A2(n2866), .ZN(n3070) );
  OAI22_X1 U2560 ( .A1(n949), .A2(n3071), .B1(n3072), .B2(n3073), .ZN(n1111)
         );
  INV_X1 U2561 ( .A(sum[0]), .ZN(n3072) );
  OAI22_X1 U2562 ( .A1(n948), .A2(n3071), .B1(n3074), .B2(n3073), .ZN(n1110)
         );
  INV_X1 U2563 ( .A(sum[1]), .ZN(n3074) );
  OAI22_X1 U2564 ( .A1(n947), .A2(n3071), .B1(n3075), .B2(n3073), .ZN(n1109)
         );
  INV_X1 U2565 ( .A(sum[2]), .ZN(n3075) );
  OAI22_X1 U2566 ( .A1(n946), .A2(n3071), .B1(n3076), .B2(n3073), .ZN(n1108)
         );
  INV_X1 U2567 ( .A(sum[3]), .ZN(n3076) );
  OAI22_X1 U2568 ( .A1(n945), .A2(n3071), .B1(n3077), .B2(n3073), .ZN(n1107)
         );
  INV_X1 U2569 ( .A(sum[4]), .ZN(n3077) );
  OAI22_X1 U2570 ( .A1(n944), .A2(n3071), .B1(n3078), .B2(n3073), .ZN(n1106)
         );
  NAND2_X1 U2571 ( .A1(n3079), .A2(n3071), .ZN(n3073) );
  INV_X1 U2572 ( .A(n2876), .ZN(n3079) );
  INV_X1 U2573 ( .A(sum[5]), .ZN(n3078) );
  OAI21_X1 U2574 ( .B1(n3305), .B2(n2876), .A(n2985), .ZN(n3071) );
  MUX2_X1 U2575 ( .A(nq[0]), .B(n3080), .S(n3081), .Z(n1105) );
  MUX2_X1 U2576 ( .A(nq[1]), .B(n3080), .S(n3082), .Z(n1104) );
  MUX2_X1 U2577 ( .A(nq[2]), .B(n3080), .S(n3083), .Z(n1103) );
  MUX2_X1 U2578 ( .A(nq[3]), .B(n3080), .S(n3084), .Z(n1102) );
  MUX2_X1 U2579 ( .A(nq[4]), .B(n3080), .S(n3085), .Z(n1101) );
  MUX2_X1 U2580 ( .A(nq[5]), .B(n3080), .S(n3086), .Z(n1100) );
  MUX2_X1 U2581 ( .A(nq[6]), .B(n3080), .S(n3087), .Z(n1099) );
  MUX2_X1 U2582 ( .A(nq[7]), .B(n3080), .S(n3088), .Z(n1098) );
  MUX2_X1 U2583 ( .A(nq[8]), .B(n3080), .S(n3089), .Z(n1097) );
  MUX2_X1 U2584 ( .A(nq[9]), .B(n3080), .S(n3090), .Z(n1096) );
  MUX2_X1 U2585 ( .A(nq[10]), .B(n3080), .S(n3091), .Z(n1095) );
  MUX2_X1 U2586 ( .A(nq[11]), .B(n3080), .S(n3092), .Z(n1094) );
  MUX2_X1 U2587 ( .A(nq[12]), .B(n3080), .S(n3093), .Z(n1093) );
  MUX2_X1 U2588 ( .A(nq[13]), .B(n3080), .S(n3094), .Z(n1092) );
  MUX2_X1 U2589 ( .A(nq[14]), .B(n3080), .S(n3095), .Z(n1091) );
  MUX2_X1 U2590 ( .A(nq[15]), .B(n3080), .S(n3096), .Z(n1090) );
  MUX2_X1 U2591 ( .A(nq[16]), .B(n3080), .S(n3097), .Z(n1089) );
  MUX2_X1 U2592 ( .A(nq[17]), .B(n3080), .S(n3098), .Z(n1088) );
  MUX2_X1 U2593 ( .A(nq[18]), .B(n3080), .S(n3099), .Z(n1087) );
  MUX2_X1 U2594 ( .A(nq[19]), .B(n3080), .S(n3100), .Z(n1086) );
  MUX2_X1 U2595 ( .A(nq[20]), .B(n3080), .S(n3101), .Z(n1085) );
  MUX2_X1 U2596 ( .A(nq[21]), .B(n3080), .S(n3102), .Z(n1084) );
  MUX2_X1 U2597 ( .A(nq[22]), .B(n3080), .S(n3103), .Z(n1083) );
  MUX2_X1 U2598 ( .A(nq[23]), .B(n3080), .S(n3104), .Z(n1082) );
  MUX2_X1 U2599 ( .A(nq[24]), .B(n3080), .S(n3105), .Z(n1081) );
  MUX2_X1 U2600 ( .A(nq[25]), .B(n3080), .S(n3106), .Z(n1080) );
  MUX2_X1 U2601 ( .A(nq[26]), .B(n3080), .S(n3107), .Z(n1079) );
  MUX2_X1 U2602 ( .A(nq[27]), .B(n3080), .S(n3108), .Z(n1078) );
  MUX2_X1 U2603 ( .A(nq[28]), .B(n3080), .S(n3109), .Z(n1077) );
  MUX2_X1 U2604 ( .A(nq[29]), .B(n3080), .S(n3110), .Z(n1076) );
  MUX2_X1 U2605 ( .A(nq[30]), .B(n3080), .S(n3111), .Z(n1075) );
  MUX2_X1 U2606 ( .A(q[0]), .B(n3113), .S(n3081), .Z(n1074) );
  OAI21_X1 U2607 ( .B1(n3114), .B2(n3115), .A(n2995), .ZN(n3081) );
  MUX2_X1 U2608 ( .A(q[1]), .B(n3113), .S(n3082), .Z(n1073) );
  OAI21_X1 U2609 ( .B1(n3114), .B2(n3116), .A(n2995), .ZN(n3082) );
  MUX2_X1 U2610 ( .A(q[2]), .B(n3113), .S(n3083), .Z(n1072) );
  OAI21_X1 U2611 ( .B1(n3114), .B2(n3117), .A(n2995), .ZN(n3083) );
  MUX2_X1 U2612 ( .A(q[3]), .B(n3113), .S(n3084), .Z(n1071) );
  OAI21_X1 U2613 ( .B1(n3114), .B2(n3118), .A(n2995), .ZN(n3084) );
  MUX2_X1 U2614 ( .A(q[4]), .B(n3113), .S(n3085), .Z(n1070) );
  OAI21_X1 U2615 ( .B1(n3114), .B2(n3119), .A(n2995), .ZN(n3085) );
  MUX2_X1 U2616 ( .A(q[5]), .B(n3113), .S(n3086), .Z(n1069) );
  OAI21_X1 U2617 ( .B1(n3114), .B2(n3120), .A(n2995), .ZN(n3086) );
  MUX2_X1 U2618 ( .A(q[6]), .B(n3113), .S(n3087), .Z(n1068) );
  OAI21_X1 U2619 ( .B1(n3114), .B2(n3121), .A(n2995), .ZN(n3087) );
  MUX2_X1 U2620 ( .A(q[7]), .B(n3113), .S(n3088), .Z(n1067) );
  OAI21_X1 U2621 ( .B1(n3114), .B2(n3122), .A(n2995), .ZN(n3088) );
  NAND3_X1 U2622 ( .A1(n935), .A2(n2929), .A3(n936), .ZN(n3114) );
  MUX2_X1 U2623 ( .A(q[8]), .B(n3113), .S(n3089), .Z(n1066) );
  OAI21_X1 U2624 ( .B1(n3115), .B2(n3123), .A(n2995), .ZN(n3089) );
  MUX2_X1 U2625 ( .A(q[9]), .B(n3113), .S(n3090), .Z(n1065) );
  OAI21_X1 U2626 ( .B1(n3116), .B2(n3123), .A(n2995), .ZN(n3090) );
  MUX2_X1 U2627 ( .A(q[10]), .B(n3113), .S(n3091), .Z(n1064) );
  OAI21_X1 U2628 ( .B1(n3117), .B2(n3123), .A(n2995), .ZN(n3091) );
  MUX2_X1 U2629 ( .A(q[11]), .B(n3113), .S(n3092), .Z(n1063) );
  OAI21_X1 U2630 ( .B1(n3118), .B2(n3123), .A(n2995), .ZN(n3092) );
  MUX2_X1 U2631 ( .A(q[12]), .B(n3113), .S(n3093), .Z(n1062) );
  OAI21_X1 U2632 ( .B1(n3119), .B2(n3123), .A(n2995), .ZN(n3093) );
  MUX2_X1 U2633 ( .A(q[13]), .B(n3113), .S(n3094), .Z(n1061) );
  OAI21_X1 U2634 ( .B1(n3120), .B2(n3123), .A(n2995), .ZN(n3094) );
  MUX2_X1 U2635 ( .A(q[14]), .B(n3113), .S(n3095), .Z(n1060) );
  OAI21_X1 U2636 ( .B1(n3121), .B2(n3123), .A(n2995), .ZN(n3095) );
  MUX2_X1 U2637 ( .A(q[15]), .B(n3113), .S(n3096), .Z(n1059) );
  OAI21_X1 U2638 ( .B1(n3122), .B2(n3123), .A(n2995), .ZN(n3096) );
  NAND3_X1 U2639 ( .A1(n2929), .A2(ct[3]), .A3(n935), .ZN(n3123) );
  MUX2_X1 U2640 ( .A(q[16]), .B(n3113), .S(n3097), .Z(n1058) );
  OAI21_X1 U2641 ( .B1(n3115), .B2(n3124), .A(n2995), .ZN(n3097) );
  MUX2_X1 U2642 ( .A(q[17]), .B(n3113), .S(n3098), .Z(n1057) );
  OAI21_X1 U2643 ( .B1(n3116), .B2(n3124), .A(n2995), .ZN(n3098) );
  MUX2_X1 U2644 ( .A(q[18]), .B(n3113), .S(n3099), .Z(n1056) );
  OAI21_X1 U2645 ( .B1(n3117), .B2(n3124), .A(n2995), .ZN(n3099) );
  MUX2_X1 U2646 ( .A(q[19]), .B(n3113), .S(n3100), .Z(n1055) );
  OAI21_X1 U2647 ( .B1(n3118), .B2(n3124), .A(n2995), .ZN(n3100) );
  MUX2_X1 U2648 ( .A(q[20]), .B(n3113), .S(n3101), .Z(n1054) );
  OAI21_X1 U2649 ( .B1(n3119), .B2(n3124), .A(n2995), .ZN(n3101) );
  MUX2_X1 U2650 ( .A(q[21]), .B(n3113), .S(n3102), .Z(n1053) );
  OAI21_X1 U2651 ( .B1(n3120), .B2(n3124), .A(n2995), .ZN(n3102) );
  MUX2_X1 U2652 ( .A(q[22]), .B(n3113), .S(n3103), .Z(n1052) );
  OAI21_X1 U2653 ( .B1(n3121), .B2(n3124), .A(n2995), .ZN(n3103) );
  MUX2_X1 U2654 ( .A(q[23]), .B(n3113), .S(n3104), .Z(n1051) );
  OAI21_X1 U2655 ( .B1(n3122), .B2(n3124), .A(n2995), .ZN(n3104) );
  NAND3_X1 U2656 ( .A1(n2929), .A2(ct[4]), .A3(n936), .ZN(n3124) );
  NAND3_X1 U2657 ( .A1(ct[1]), .A2(ct[0]), .A3(ct[2]), .ZN(n3122) );
  MUX2_X1 U2658 ( .A(q[24]), .B(n3113), .S(n3105), .Z(n1050) );
  OAI21_X1 U2659 ( .B1(n3115), .B2(n3125), .A(n2995), .ZN(n3105) );
  NAND3_X1 U2660 ( .A1(n938), .A2(n937), .A3(n939), .ZN(n3115) );
  MUX2_X1 U2661 ( .A(q[25]), .B(n3113), .S(n3106), .Z(n1049) );
  OAI21_X1 U2662 ( .B1(n3116), .B2(n3125), .A(n2995), .ZN(n3106) );
  NAND3_X1 U2663 ( .A1(n937), .A2(ct[0]), .A3(n938), .ZN(n3116) );
  MUX2_X1 U2664 ( .A(q[26]), .B(n3113), .S(n3107), .Z(n1048) );
  OAI21_X1 U2665 ( .B1(n3117), .B2(n3125), .A(n2995), .ZN(n3107) );
  NAND3_X1 U2666 ( .A1(n937), .A2(ct[1]), .A3(n939), .ZN(n3117) );
  MUX2_X1 U2667 ( .A(q[27]), .B(n3113), .S(n3108), .Z(n1047) );
  OAI21_X1 U2668 ( .B1(n3118), .B2(n3125), .A(n2995), .ZN(n3108) );
  NAND3_X1 U2669 ( .A1(ct[1]), .A2(ct[0]), .A3(n937), .ZN(n3118) );
  MUX2_X1 U2670 ( .A(q[28]), .B(n3113), .S(n3109), .Z(n1046) );
  OAI21_X1 U2671 ( .B1(n3119), .B2(n3125), .A(n2995), .ZN(n3109) );
  NAND3_X1 U2672 ( .A1(n938), .A2(ct[2]), .A3(n939), .ZN(n3119) );
  MUX2_X1 U2673 ( .A(q[29]), .B(n3113), .S(n3110), .Z(n1045) );
  OAI21_X1 U2674 ( .B1(n3120), .B2(n3125), .A(n2995), .ZN(n3110) );
  NAND3_X1 U2675 ( .A1(ct[2]), .A2(ct[0]), .A3(n938), .ZN(n3120) );
  MUX2_X1 U2676 ( .A(q[30]), .B(n3113), .S(n3111), .Z(n1044) );
  OAI21_X1 U2677 ( .B1(n3121), .B2(n3125), .A(n2995), .ZN(n3111) );
  AND4_X1 U2678 ( .A1(state[0]), .A2(n3126), .A3(n2799), .A4(n2855), .ZN(n2986) );
  NAND3_X1 U2679 ( .A1(ct[4]), .A2(ct[3]), .A3(n2929), .ZN(n3125) );
  INV_X1 U2680 ( .A(n2943), .ZN(n2929) );
  NAND3_X1 U2681 ( .A1(n2991), .A2(n2998), .A3(n934), .ZN(n2943) );
  INV_X1 U2682 ( .A(n2878), .ZN(n2991) );
  NAND3_X1 U2683 ( .A1(ct[2]), .A2(ct[1]), .A3(n939), .ZN(n3121) );
  NAND4_X1 U2684 ( .A1(state[2]), .A2(n3126), .A3(n2807), .A4(n2799), .ZN(
        n2878) );
  OAI221_X1 U2685 ( .B1(n3128), .B2(n3129), .C1(n2927), .C2(n940), .A(n2982), 
        .ZN(n1043) );
  AOI21_X1 U2686 ( .B1(n3112), .B2(n3130), .A(n2983), .ZN(n3128) );
  INV_X1 U2687 ( .A(n2984), .ZN(n2983) );
  OR4_X1 U2688 ( .A1(n3131), .A2(n3132), .A3(n3133), .A4(n3134), .ZN(n1042) );
  OAI222_X1 U2689 ( .A1(nqp1[0]), .A2(n3135), .B1(n3301), .B2(n2933), .C1(
        nq[0]), .C2(n3136), .ZN(n3134) );
  MUX2_X1 U2690 ( .A(n2861), .B(n2859), .S(i_divisor[0]), .Z(n3133) );
  MUX2_X1 U2691 ( .A(n3137), .B(n2860), .S(n3306), .Z(n3132) );
  NOR2_X1 U2692 ( .A1(n2927), .A2(n1773), .ZN(n3131) );
  OR4_X1 U2693 ( .A1(n3138), .A2(n3139), .A3(n3140), .A4(n3141), .ZN(n1041) );
  OAI222_X1 U2694 ( .A1(nqp1[1]), .A2(n3135), .B1(n3302), .B2(n2933), .C1(
        nq[1]), .C2(n3136), .ZN(n3141) );
  MUX2_X1 U2695 ( .A(n2861), .B(n2859), .S(i_divisor[1]), .Z(n3140) );
  MUX2_X1 U2696 ( .A(n3137), .B(n2860), .S(n3341), .Z(n3139) );
  NOR2_X1 U2697 ( .A1(n2927), .A2(n1772), .ZN(n3138) );
  OR4_X1 U2698 ( .A1(n3142), .A2(n3143), .A3(n3144), .A4(n3145), .ZN(n1040) );
  OAI222_X1 U2699 ( .A1(nqp1[2]), .A2(n3135), .B1(n3303), .B2(n2933), .C1(
        nq[2]), .C2(n3136), .ZN(n3145) );
  MUX2_X1 U2700 ( .A(n2861), .B(n2859), .S(i_divisor[2]), .Z(n3144) );
  MUX2_X1 U2701 ( .A(n3137), .B(n2860), .S(n3339), .Z(n3143) );
  NOR2_X1 U2702 ( .A1(n2927), .A2(n1771), .ZN(n3142) );
  OR4_X1 U2703 ( .A1(n3146), .A2(n3147), .A3(n3148), .A4(n3149), .ZN(n1039) );
  OAI222_X1 U2704 ( .A1(nqp1[3]), .A2(n3135), .B1(n3304), .B2(n2933), .C1(
        nq[3]), .C2(n3136), .ZN(n3149) );
  MUX2_X1 U2705 ( .A(n2861), .B(n2859), .S(i_divisor[3]), .Z(n3148) );
  MUX2_X1 U2706 ( .A(n3137), .B(n2860), .S(n3337), .Z(n3147) );
  NOR2_X1 U2707 ( .A1(n2927), .A2(n1770), .ZN(n3146) );
  OR4_X1 U2708 ( .A1(n3150), .A2(n3151), .A3(n3152), .A4(n3153), .ZN(n1038) );
  NAND2_X1 U2709 ( .A1(n3298), .A2(n2927), .ZN(n2933) );
  MUX2_X1 U2710 ( .A(n2861), .B(n2859), .S(i_divisor[4]), .Z(n3152) );
  MUX2_X1 U2711 ( .A(n3137), .B(n2860), .S(n3335), .Z(n3151) );
  NOR2_X1 U2712 ( .A1(n2927), .A2(n1769), .ZN(n3150) );
  OR3_X1 U2713 ( .A1(n3154), .A2(n3155), .A3(n3156), .ZN(n1037) );
  OAI222_X1 U2714 ( .A1(nq[5]), .A2(n3136), .B1(nqp1[5]), .B2(n3135), .C1(
        n2927), .C2(n802), .ZN(n3156) );
  MUX2_X1 U2715 ( .A(n3137), .B(n2860), .S(n3333), .Z(n3155) );
  MUX2_X1 U2716 ( .A(n2861), .B(n2859), .S(i_divisor[5]), .Z(n3154) );
  OR3_X1 U2717 ( .A1(n3157), .A2(n3158), .A3(n3159), .ZN(n1036) );
  OAI222_X1 U2718 ( .A1(nq[6]), .A2(n3136), .B1(nqp1[6]), .B2(n3135), .C1(
        n2927), .C2(n803), .ZN(n3159) );
  MUX2_X1 U2719 ( .A(n3137), .B(n2860), .S(n3332), .Z(n3158) );
  MUX2_X1 U2720 ( .A(n2861), .B(n2859), .S(i_divisor[6]), .Z(n3157) );
  OR3_X1 U2721 ( .A1(n3160), .A2(n3161), .A3(n3162), .ZN(n1035) );
  OAI222_X1 U2722 ( .A1(nq[7]), .A2(n3136), .B1(nqp1[7]), .B2(n3135), .C1(
        n2927), .C2(n804), .ZN(n3162) );
  MUX2_X1 U2723 ( .A(n3137), .B(n2860), .S(n3331), .Z(n3161) );
  MUX2_X1 U2724 ( .A(n2861), .B(n2859), .S(i_divisor[7]), .Z(n3160) );
  OR3_X1 U2725 ( .A1(n3163), .A2(n3164), .A3(n3165), .ZN(n1034) );
  OAI222_X1 U2726 ( .A1(nq[8]), .A2(n3136), .B1(nqp1[8]), .B2(n3135), .C1(
        n2927), .C2(n805), .ZN(n3165) );
  MUX2_X1 U2727 ( .A(n3137), .B(n2860), .S(n3330), .Z(n3164) );
  MUX2_X1 U2728 ( .A(n2861), .B(n2859), .S(i_divisor[8]), .Z(n3163) );
  OR3_X1 U2729 ( .A1(n3166), .A2(n3167), .A3(n3168), .ZN(n1033) );
  OAI222_X1 U2730 ( .A1(nq[9]), .A2(n3136), .B1(nqp1[9]), .B2(n3135), .C1(
        n2927), .C2(n806), .ZN(n3168) );
  MUX2_X1 U2731 ( .A(n3137), .B(n2860), .S(n3329), .Z(n3167) );
  MUX2_X1 U2732 ( .A(n2861), .B(n2859), .S(i_divisor[9]), .Z(n3166) );
  OR3_X1 U2733 ( .A1(n3169), .A2(n3170), .A3(n3171), .ZN(n1032) );
  OAI222_X1 U2734 ( .A1(nq[10]), .A2(n3136), .B1(nqp1[10]), .B2(n3135), .C1(
        n2927), .C2(n807), .ZN(n3171) );
  MUX2_X1 U2735 ( .A(n3137), .B(n2860), .S(n3328), .Z(n3170) );
  MUX2_X1 U2736 ( .A(n2861), .B(n2859), .S(i_divisor[10]), .Z(n3169) );
  OR3_X1 U2737 ( .A1(n3172), .A2(n3173), .A3(n3174), .ZN(n1031) );
  OAI222_X1 U2738 ( .A1(nq[11]), .A2(n3136), .B1(nqp1[11]), .B2(n3135), .C1(
        n2927), .C2(n808), .ZN(n3174) );
  MUX2_X1 U2739 ( .A(n3137), .B(n2860), .S(n3327), .Z(n3173) );
  MUX2_X1 U2740 ( .A(n2861), .B(n2859), .S(i_divisor[11]), .Z(n3172) );
  OR3_X1 U2741 ( .A1(n3175), .A2(n3176), .A3(n3177), .ZN(n1030) );
  OAI222_X1 U2742 ( .A1(nq[12]), .A2(n3136), .B1(nqp1[12]), .B2(n3135), .C1(
        n2927), .C2(n809), .ZN(n3177) );
  MUX2_X1 U2743 ( .A(n3137), .B(n2860), .S(n3326), .Z(n3176) );
  MUX2_X1 U2744 ( .A(n2861), .B(n2859), .S(i_divisor[12]), .Z(n3175) );
  OR3_X1 U2745 ( .A1(n3178), .A2(n3179), .A3(n3180), .ZN(n1029) );
  OAI222_X1 U2746 ( .A1(nq[13]), .A2(n3136), .B1(nqp1[13]), .B2(n3135), .C1(
        n2927), .C2(n810), .ZN(n3180) );
  MUX2_X1 U2747 ( .A(n3137), .B(n2860), .S(n3325), .Z(n3179) );
  MUX2_X1 U2748 ( .A(n2861), .B(n2859), .S(i_divisor[13]), .Z(n3178) );
  OR3_X1 U2749 ( .A1(n3181), .A2(n3182), .A3(n3183), .ZN(n1028) );
  OAI222_X1 U2750 ( .A1(nq[14]), .A2(n3136), .B1(nqp1[14]), .B2(n3135), .C1(
        n2927), .C2(n811), .ZN(n3183) );
  MUX2_X1 U2751 ( .A(n3137), .B(n2860), .S(n3324), .Z(n3182) );
  MUX2_X1 U2752 ( .A(n2861), .B(n2859), .S(i_divisor[14]), .Z(n3181) );
  OR3_X1 U2753 ( .A1(n3184), .A2(n3185), .A3(n3186), .ZN(n1027) );
  OAI222_X1 U2754 ( .A1(nq[15]), .A2(n3136), .B1(nqp1[15]), .B2(n3135), .C1(
        n2927), .C2(n812), .ZN(n3186) );
  MUX2_X1 U2755 ( .A(n3137), .B(n2860), .S(n3323), .Z(n3185) );
  MUX2_X1 U2756 ( .A(n2861), .B(n2859), .S(i_divisor[15]), .Z(n3184) );
  OR3_X1 U2757 ( .A1(n3187), .A2(n3188), .A3(n3189), .ZN(n1026) );
  OAI222_X1 U2758 ( .A1(nq[16]), .A2(n3136), .B1(nqp1[16]), .B2(n3135), .C1(
        n2927), .C2(n813), .ZN(n3189) );
  MUX2_X1 U2759 ( .A(n3137), .B(n2860), .S(n3322), .Z(n3188) );
  MUX2_X1 U2760 ( .A(n2861), .B(n2859), .S(i_divisor[16]), .Z(n3187) );
  OR3_X1 U2761 ( .A1(n3190), .A2(n3191), .A3(n3192), .ZN(n1025) );
  OAI222_X1 U2762 ( .A1(nq[17]), .A2(n3136), .B1(nqp1[17]), .B2(n3135), .C1(
        n2927), .C2(n814), .ZN(n3192) );
  MUX2_X1 U2763 ( .A(n3137), .B(n2860), .S(n3321), .Z(n3191) );
  MUX2_X1 U2764 ( .A(n2861), .B(n2859), .S(i_divisor[17]), .Z(n3190) );
  OR3_X1 U2765 ( .A1(n3193), .A2(n3194), .A3(n3195), .ZN(n1024) );
  OAI222_X1 U2766 ( .A1(nq[18]), .A2(n3136), .B1(nqp1[18]), .B2(n3135), .C1(
        n2927), .C2(n815), .ZN(n3195) );
  MUX2_X1 U2767 ( .A(n3137), .B(n2860), .S(n3320), .Z(n3194) );
  MUX2_X1 U2768 ( .A(n2861), .B(n2859), .S(i_divisor[18]), .Z(n3193) );
  OR3_X1 U2769 ( .A1(n3196), .A2(n3197), .A3(n3198), .ZN(n1023) );
  OAI222_X1 U2770 ( .A1(nq[19]), .A2(n3136), .B1(nqp1[19]), .B2(n3135), .C1(
        n2927), .C2(n816), .ZN(n3198) );
  MUX2_X1 U2771 ( .A(n3137), .B(n2860), .S(n3319), .Z(n3197) );
  MUX2_X1 U2772 ( .A(n2861), .B(n2859), .S(i_divisor[19]), .Z(n3196) );
  OR3_X1 U2773 ( .A1(n3199), .A2(n3200), .A3(n3201), .ZN(n1022) );
  OAI222_X1 U2774 ( .A1(nq[20]), .A2(n3136), .B1(nqp1[20]), .B2(n3135), .C1(
        n2927), .C2(n817), .ZN(n3201) );
  MUX2_X1 U2775 ( .A(n3137), .B(n2860), .S(n3318), .Z(n3200) );
  MUX2_X1 U2776 ( .A(n2861), .B(n2859), .S(i_divisor[20]), .Z(n3199) );
  OR3_X1 U2777 ( .A1(n3202), .A2(n3203), .A3(n3204), .ZN(n1021) );
  OAI222_X1 U2778 ( .A1(nq[21]), .A2(n3136), .B1(nqp1[21]), .B2(n3135), .C1(
        n2927), .C2(n818), .ZN(n3204) );
  MUX2_X1 U2779 ( .A(n3137), .B(n2860), .S(n3317), .Z(n3203) );
  MUX2_X1 U2780 ( .A(n2861), .B(n2859), .S(i_divisor[21]), .Z(n3202) );
  OR3_X1 U2781 ( .A1(n3205), .A2(n3206), .A3(n3207), .ZN(n1020) );
  OAI222_X1 U2782 ( .A1(nq[22]), .A2(n3136), .B1(nqp1[22]), .B2(n3135), .C1(
        n2927), .C2(n819), .ZN(n3207) );
  MUX2_X1 U2783 ( .A(n3137), .B(n2860), .S(n3316), .Z(n3206) );
  MUX2_X1 U2784 ( .A(n2861), .B(n2859), .S(i_divisor[22]), .Z(n3205) );
  OR3_X1 U2785 ( .A1(n3208), .A2(n3209), .A3(n3210), .ZN(n1019) );
  OAI222_X1 U2786 ( .A1(nq[23]), .A2(n3136), .B1(nqp1[23]), .B2(n3135), .C1(
        n2927), .C2(n820), .ZN(n3210) );
  MUX2_X1 U2787 ( .A(n3137), .B(n2860), .S(n3315), .Z(n3209) );
  MUX2_X1 U2788 ( .A(n2861), .B(n2859), .S(i_divisor[23]), .Z(n3208) );
  OR3_X1 U2789 ( .A1(n3211), .A2(n3212), .A3(n3213), .ZN(n1018) );
  OAI222_X1 U2790 ( .A1(nq[24]), .A2(n3136), .B1(nqp1[24]), .B2(n3135), .C1(
        n2927), .C2(n821), .ZN(n3213) );
  MUX2_X1 U2791 ( .A(n3137), .B(n2860), .S(n3314), .Z(n3212) );
  MUX2_X1 U2792 ( .A(n2861), .B(n2859), .S(i_divisor[24]), .Z(n3211) );
  OR3_X1 U2793 ( .A1(n3214), .A2(n3215), .A3(n3216), .ZN(n1017) );
  OAI222_X1 U2794 ( .A1(nq[25]), .A2(n3136), .B1(nqp1[25]), .B2(n3135), .C1(
        n2927), .C2(n822), .ZN(n3216) );
  MUX2_X1 U2795 ( .A(n3137), .B(n2860), .S(n3313), .Z(n3215) );
  MUX2_X1 U2796 ( .A(n2861), .B(n2859), .S(i_divisor[25]), .Z(n3214) );
  OR3_X1 U2797 ( .A1(n3217), .A2(n3218), .A3(n3219), .ZN(n1016) );
  OAI222_X1 U2798 ( .A1(nq[26]), .A2(n3136), .B1(nqp1[26]), .B2(n3135), .C1(
        n2927), .C2(n823), .ZN(n3219) );
  MUX2_X1 U2799 ( .A(n3137), .B(n2860), .S(n3312), .Z(n3218) );
  MUX2_X1 U2800 ( .A(n2861), .B(n2859), .S(i_divisor[26]), .Z(n3217) );
  OR3_X1 U2801 ( .A1(n3220), .A2(n3221), .A3(n3222), .ZN(n1015) );
  OAI222_X1 U2802 ( .A1(nq[27]), .A2(n3136), .B1(nqp1[27]), .B2(n3135), .C1(
        n2927), .C2(n824), .ZN(n3222) );
  MUX2_X1 U2803 ( .A(n3137), .B(n2860), .S(n3311), .Z(n3221) );
  MUX2_X1 U2804 ( .A(n2861), .B(n2859), .S(i_divisor[27]), .Z(n3220) );
  OR3_X1 U2805 ( .A1(n3223), .A2(n3224), .A3(n3225), .ZN(n1014) );
  OAI222_X1 U2806 ( .A1(nq[28]), .A2(n3136), .B1(nqp1[28]), .B2(n3135), .C1(
        n2927), .C2(n825), .ZN(n3225) );
  MUX2_X1 U2807 ( .A(n3137), .B(n2860), .S(n3310), .Z(n3224) );
  MUX2_X1 U2808 ( .A(n2861), .B(n2859), .S(i_divisor[28]), .Z(n3223) );
  OR3_X1 U2809 ( .A1(n3226), .A2(n3227), .A3(n3228), .ZN(n1013) );
  OAI222_X1 U2810 ( .A1(nq[29]), .A2(n3136), .B1(nqp1[29]), .B2(n3135), .C1(
        n2927), .C2(n826), .ZN(n3228) );
  MUX2_X1 U2811 ( .A(n3137), .B(n2860), .S(n3309), .Z(n3227) );
  MUX2_X1 U2812 ( .A(n2861), .B(n2859), .S(i_divisor[29]), .Z(n3226) );
  OR3_X1 U2813 ( .A1(n3229), .A2(n3230), .A3(n3231), .ZN(n1012) );
  OAI222_X1 U2814 ( .A1(nq[30]), .A2(n3136), .B1(nqp1[30]), .B2(n3135), .C1(
        n2927), .C2(n827), .ZN(n3231) );
  MUX2_X1 U2815 ( .A(n3137), .B(n2860), .S(n3308), .Z(n3230) );
  MUX2_X1 U2816 ( .A(n2861), .B(n2859), .S(i_divisor[30]), .Z(n3229) );
  OR3_X1 U2817 ( .A1(n3234), .A2(n3235), .A3(n3236), .ZN(n1011) );
  OAI21_X1 U2818 ( .B1(n2857), .B2(n2927), .A(n2982), .ZN(n3236) );
  INV_X1 U2819 ( .A(n3233), .ZN(n2982) );
  NOR2_X1 U2820 ( .A1(n3129), .A2(n3237), .ZN(n3233) );
  MUX2_X1 U2821 ( .A(n2861), .B(n2859), .S(i_divisor[31]), .Z(n3235) );
  NAND2_X1 U2822 ( .A1(n3127), .A2(n3238), .ZN(n3232) );
  INV_X1 U2823 ( .A(n2935), .ZN(n2926) );
  NAND2_X1 U2824 ( .A1(n3238), .A2(n3112), .ZN(n2984) );
  MUX2_X1 U2825 ( .A(n2854), .B(n3239), .S(n3307), .Z(n3238) );
  AOI21_X1 U2826 ( .B1(n3240), .B2(n3241), .A(n2854), .ZN(n3239) );
  NOR4_X1 U2827 ( .A1(n3242), .A2(n3243), .A3(n3244), .A4(n3245), .ZN(n3241)
         );
  NAND4_X1 U2828 ( .A1(n2847), .A2(n2800), .A3(n2793), .A4(n2787), .ZN(n3245)
         );
  NAND4_X1 U2829 ( .A1(n2848), .A2(n2801), .A3(n2794), .A4(n2788), .ZN(n3244)
         );
  NAND4_X1 U2830 ( .A1(n2849), .A2(n2802), .A3(n2795), .A4(n2789), .ZN(n3243)
         );
  NAND4_X1 U2831 ( .A1(n2850), .A2(n2803), .A3(n2796), .A4(n2790), .ZN(n3242)
         );
  NOR4_X1 U2832 ( .A1(n3246), .A2(n3247), .A3(n3248), .A4(n3249), .ZN(n3240)
         );
  OR3_X1 U2833 ( .A1(n3342), .A2(n3340), .A3(n3348), .ZN(n3249) );
  OR4_X1 U2834 ( .A1(n3338), .A2(n3336), .A3(n3334), .A4(n3297), .ZN(n3248) );
  NAND4_X1 U2835 ( .A1(n2851), .A2(n2804), .A3(n2797), .A4(n2791), .ZN(n3247)
         );
  NAND4_X1 U2836 ( .A1(n2852), .A2(n2805), .A3(n2798), .A4(n2792), .ZN(n3246)
         );
  MUX2_X1 U2837 ( .A(n3137), .B(n2860), .S(n3299), .Z(n3234) );
  INV_X1 U2838 ( .A(n3112), .ZN(n3127) );
  XOR2_X1 U2839 ( .A(n3299), .B(n3307), .Z(n3112) );
  NOR3_X1 U2840 ( .A1(n2993), .A2(n2992), .A3(n3129), .ZN(n2947) );
  OR2_X1 U2841 ( .A1(n2946), .A2(n3298), .ZN(n3129) );
  INV_X1 U2842 ( .A(n2927), .ZN(n2946) );
  NAND2_X1 U2843 ( .A1(state_reg_1_0), .A2(n941), .ZN(n2876) );
  INV_X1 U2844 ( .A(n3130), .ZN(n2993) );
  NAND4_X1 U2845 ( .A1(state[4]), .A2(n3069), .A3(n2853), .A4(n1988), .ZN(
        n3130) );
  OAI221_X1 U2846 ( .B1(n2880), .B2(n2825), .C1(n2881), .C2(n3250), .A(n3251), 
        .ZN(n1010) );
  AOI22_X1 U2847 ( .A1(n2864), .A2(PR_1[0]), .B1(N264), .B2(n2884), .ZN(n3251)
         );
  INV_X1 U2848 ( .A(i_dividend[0]), .ZN(n3250) );
  OAI221_X1 U2849 ( .B1(n2880), .B2(n2826), .C1(n2881), .C2(n3252), .A(n3253), 
        .ZN(n1009) );
  AOI22_X1 U2850 ( .A1(n2864), .A2(PR_1[1]), .B1(N265), .B2(n2884), .ZN(n3253)
         );
  INV_X1 U2851 ( .A(i_dividend[1]), .ZN(n3252) );
  OAI221_X1 U2852 ( .B1(n2880), .B2(n2827), .C1(n2881), .C2(n3254), .A(n3255), 
        .ZN(n1008) );
  AOI22_X1 U2853 ( .A1(n2864), .A2(PR_1[2]), .B1(N266), .B2(n2884), .ZN(n3255)
         );
  INV_X1 U2854 ( .A(i_dividend[2]), .ZN(n3254) );
  OAI221_X1 U2855 ( .B1(n2880), .B2(n2828), .C1(n2881), .C2(n3256), .A(n3257), 
        .ZN(n1007) );
  AOI22_X1 U2856 ( .A1(n2864), .A2(PR_1[3]), .B1(N267), .B2(n2884), .ZN(n3257)
         );
  INV_X1 U2857 ( .A(i_dividend[3]), .ZN(n3256) );
  OAI221_X1 U2858 ( .B1(n2880), .B2(n2829), .C1(n2881), .C2(n3258), .A(n3259), 
        .ZN(n1006) );
  AOI22_X1 U2859 ( .A1(n2864), .A2(PR_1[4]), .B1(N268), .B2(n2884), .ZN(n3259)
         );
  INV_X1 U2860 ( .A(i_dividend[4]), .ZN(n3258) );
  OAI221_X1 U2861 ( .B1(n2880), .B2(n2830), .C1(n2881), .C2(n3260), .A(n3261), 
        .ZN(n1005) );
  AOI22_X1 U2862 ( .A1(n2864), .A2(PR_1[5]), .B1(N269), .B2(n2884), .ZN(n3261)
         );
  INV_X1 U2863 ( .A(i_dividend[5]), .ZN(n3260) );
  OAI221_X1 U2864 ( .B1(n2880), .B2(n2831), .C1(n2881), .C2(n3262), .A(n3263), 
        .ZN(n1004) );
  AOI22_X1 U2865 ( .A1(n2864), .A2(PR_1[6]), .B1(N270), .B2(n2884), .ZN(n3263)
         );
  INV_X1 U2866 ( .A(i_dividend[6]), .ZN(n3262) );
  OAI221_X1 U2867 ( .B1(n2880), .B2(n2832), .C1(n2881), .C2(n3264), .A(n3265), 
        .ZN(n1003) );
  AOI22_X1 U2868 ( .A1(n2864), .A2(PR_1[7]), .B1(N271), .B2(n2884), .ZN(n3265)
         );
  INV_X1 U2869 ( .A(i_dividend[7]), .ZN(n3264) );
  OAI221_X1 U2870 ( .B1(n2880), .B2(n2833), .C1(n2881), .C2(n3266), .A(n3267), 
        .ZN(n1002) );
  AOI22_X1 U2871 ( .A1(n2864), .A2(PR_1[8]), .B1(N272), .B2(n2884), .ZN(n3267)
         );
  INV_X1 U2872 ( .A(i_dividend[8]), .ZN(n3266) );
  OAI221_X1 U2873 ( .B1(n2880), .B2(n2834), .C1(n2881), .C2(n3268), .A(n3269), 
        .ZN(n1001) );
  AOI22_X1 U2874 ( .A1(n2864), .A2(PR_1[9]), .B1(N273), .B2(n2884), .ZN(n3269)
         );
  INV_X1 U2875 ( .A(i_dividend[9]), .ZN(n3268) );
  OAI221_X1 U2876 ( .B1(n2880), .B2(n2835), .C1(n2881), .C2(n3270), .A(n3271), 
        .ZN(n1000) );
  AOI22_X1 U2877 ( .A1(n2864), .A2(PR_1[10]), .B1(N274), .B2(n2884), .ZN(n3271) );
  NAND2_X1 U2878 ( .A1(n2992), .A2(n2998), .ZN(n2997) );
  INV_X1 U2879 ( .A(n3237), .ZN(n2992) );
  NAND4_X1 U2880 ( .A1(state[3]), .A2(n3069), .A3(n2806), .A4(n1988), .ZN(
        n3237) );
  NOR3_X1 U2881 ( .A1(state[1]), .A2(state[2]), .A3(state[0]), .ZN(n3069) );
  INV_X1 U2882 ( .A(n2881), .ZN(n2989) );
  INV_X1 U2883 ( .A(i_dividend[10]), .ZN(n3270) );
  NOR2_X1 U2884 ( .A1(n3347), .A2(state_reg_1_0), .ZN(n2998) );
  AND4_X1 U2885 ( .A1(state[1]), .A2(n3126), .A3(n2807), .A4(n2855), .ZN(n2990) );
  NOR3_X1 U2886 ( .A1(state[4]), .A2(state[5]), .A3(state[3]), .ZN(n3126) );
  XOR2_X1 U2887 ( .A(state[5]), .B(n3343), .Z(n_1_net__3_) );
  XOR2_X1 U2888 ( .A(state[5]), .B(n3344), .Z(n_1_net__2_) );
  XOR2_X1 U2889 ( .A(state[5]), .B(n3345), .Z(n_1_net__1_) );
  XOR2_X1 U2890 ( .A(state[5]), .B(n3346), .Z(n_1_net__0_) );
  XNOR2_X1 \shifter_0/U36  ( .A(sdata[31]), .B(sdata[24]), .ZN(\shifter_0/n46 ) );
  INV_X1 \shifter_0/U35  ( .A(sdata[31]), .ZN(\shifter_0/n42 ) );
  XNOR2_X1 \shifter_0/U34  ( .A(sdata[31]), .B(sdata[27]), .ZN(\shifter_0/n48 ) );
  XNOR2_X1 \shifter_0/U33  ( .A(sdata[31]), .B(sdata[28]), .ZN(\shifter_0/n49 ) );
  XNOR2_X1 \shifter_0/U32  ( .A(sdata[31]), .B(sdata[29]), .ZN(\shifter_0/n38 ) );
  XOR2_X1 \shifter_0/U31  ( .A(sdata[31]), .B(sdata[30]), .Z(\shifter_0/n40 )
         );
  NAND2_X1 \shifter_0/U30  ( .A1(\shifter_0/n38 ), .A2(\shifter_0/n20 ), .ZN(
        \shifter_0/n32 ) );
  INV_X1 \shifter_0/U29  ( .A(\shifter_0/n32 ), .ZN(\shifter_0/n4 ) );
  NAND2_X1 \shifter_0/U28  ( .A1(\shifter_0/n49 ), .A2(\shifter_0/n4 ), .ZN(
        \shifter_0/n39 ) );
  NAND2_X1 \shifter_0/U27  ( .A1(\shifter_0/n48 ), .A2(\shifter_0/n25 ), .ZN(
        \shifter_0/n36 ) );
  INV_X1 \shifter_0/U26  ( .A(sdata[26]), .ZN(\shifter_0/n41 ) );
  MUX2_X1 \shifter_0/U25  ( .A(sdata[31]), .B(\shifter_0/n41 ), .S(sdata[25]), 
        .Z(\shifter_0/n47 ) );
  AOI211_X1 \shifter_0/U24  ( .C1(\shifter_0/n42 ), .C2(sdata[26]), .A(
        \shifter_0/n36 ), .B(\shifter_0/n47 ), .ZN(\shifter_0/n2 ) );
  NAND2_X1 \shifter_0/U23  ( .A1(\shifter_0/n46 ), .A2(\shifter_0/n2 ), .ZN(
        \shifter_0/n33 ) );
  INV_X1 \shifter_0/U22  ( .A(\shifter_0/n33 ), .ZN(\shifter_0/n1 ) );
  XNOR2_X1 \shifter_0/U21  ( .A(sdata[31]), .B(sdata[22]), .ZN(\shifter_0/n44 ) );
  XNOR2_X1 \shifter_0/U20  ( .A(sdata[31]), .B(sdata[23]), .ZN(\shifter_0/n45 ) );
  NAND2_X1 \shifter_0/U19  ( .A1(\shifter_0/n45 ), .A2(\shifter_0/n1 ), .ZN(
        \shifter_0/n30 ) );
  INV_X1 \shifter_0/U18  ( .A(\shifter_0/n30 ), .ZN(shifted_o[3]) );
  XNOR2_X1 \shifter_0/U17  ( .A(\shifter_0/n42 ), .B(sdata[26]), .ZN(
        \shifter_0/n43 ) );
  INV_X1 \shifter_0/U16  ( .A(\shifter_0/n36 ), .ZN(\shifter_0/n3 ) );
  XNOR2_X1 \shifter_0/U15  ( .A(\shifter_0/n41 ), .B(\shifter_0/n42 ), .ZN(
        \shifter_0/n35 ) );
  INV_X1 \shifter_0/U14  ( .A(\shifter_0/n2 ), .ZN(\shifter_0/n31 ) );
  AOI21_X1 \shifter_0/U13  ( .B1(\shifter_0/n38 ), .B2(\shifter_0/n39 ), .A(
        \shifter_0/n40 ), .ZN(\shifter_0/n37 ) );
  OAI221_X1 \shifter_0/U12  ( .B1(\shifter_0/n35 ), .B2(\shifter_0/n36 ), .C1(
        \shifter_0/n21 ), .C2(\shifter_0/n31 ), .A(\shifter_0/n37 ), .ZN(
        \shifter_0/n34 ) );
  OAI21_X1 \shifter_0/U11  ( .B1(shifted_o[3]), .B2(\shifter_0/n33 ), .A(
        \shifter_0/n34 ), .ZN(shifted_o[0]) );
  OAI22_X1 \shifter_0/U10  ( .A1(\shifter_0/n3 ), .A2(\shifter_0/n32 ), .B1(
        shifted_o[3]), .B2(\shifter_0/n31 ), .ZN(shifted_o[1]) );
  MUX2_X1 \shifter_0/U9  ( .A(\shifter_0/n30 ), .B(\shifter_0/n3 ), .S(
        \shifter_0/n31 ), .Z(shifted_o[2]) );
  NOR2_X4 \shifter_0/U8  ( .A1(\shifter_0/n36 ), .A2(\shifter_0/n43 ), .ZN(
        \shifter_0/n24 ) );
  AND2_X2 \shifter_0/U7  ( .A1(\shifter_0/n44 ), .A2(shifted_o[3]), .ZN(
        \shifter_0/n21 ) );
  INV_X2 \shifter_0/U6  ( .A(\shifter_0/n39 ), .ZN(\shifter_0/n25 ) );
  INV_X2 \shifter_0/U5  ( .A(\shifter_0/n40 ), .ZN(\shifter_0/n20 ) );
  INV_X1 \shifter_0/U3  ( .A(1'b1), .ZN(\shifter_0/o_shifted[4] ) );
  INV_X1 \shifter_0/shift_1b_0/U97  ( .A(sdata[0]), .ZN(
        \shifter_0/shift_1b_0/n33 ) );
  NOR2_X1 \shifter_0/shift_1b_0/U96  ( .A1(\shifter_0/n20 ), .A2(
        \shifter_0/shift_1b_0/n33 ), .ZN(\shifter_0/data_1 [0]) );
  MUX2_X1 \shifter_0/shift_1b_0/U95  ( .A(sdata[10]), .B(sdata[9]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [10]) );
  MUX2_X1 \shifter_0/shift_1b_0/U94  ( .A(sdata[11]), .B(sdata[10]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [11]) );
  MUX2_X1 \shifter_0/shift_1b_0/U93  ( .A(sdata[12]), .B(sdata[11]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [12]) );
  MUX2_X1 \shifter_0/shift_1b_0/U92  ( .A(sdata[13]), .B(sdata[12]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [13]) );
  MUX2_X1 \shifter_0/shift_1b_0/U91  ( .A(sdata[14]), .B(sdata[13]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [14]) );
  MUX2_X1 \shifter_0/shift_1b_0/U90  ( .A(sdata[15]), .B(sdata[14]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [15]) );
  MUX2_X1 \shifter_0/shift_1b_0/U89  ( .A(sdata[16]), .B(sdata[15]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [16]) );
  MUX2_X1 \shifter_0/shift_1b_0/U88  ( .A(sdata[17]), .B(sdata[16]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [17]) );
  MUX2_X1 \shifter_0/shift_1b_0/U87  ( .A(sdata[18]), .B(sdata[17]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [18]) );
  MUX2_X1 \shifter_0/shift_1b_0/U86  ( .A(sdata[19]), .B(sdata[18]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [19]) );
  MUX2_X1 \shifter_0/shift_1b_0/U85  ( .A(sdata[1]), .B(sdata[0]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [1]) );
  MUX2_X1 \shifter_0/shift_1b_0/U84  ( .A(sdata[20]), .B(sdata[19]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [20]) );
  MUX2_X1 \shifter_0/shift_1b_0/U83  ( .A(sdata[21]), .B(sdata[20]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [21]) );
  MUX2_X1 \shifter_0/shift_1b_0/U82  ( .A(sdata[22]), .B(sdata[21]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [22]) );
  MUX2_X1 \shifter_0/shift_1b_0/U81  ( .A(sdata[23]), .B(sdata[22]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [23]) );
  MUX2_X1 \shifter_0/shift_1b_0/U80  ( .A(sdata[24]), .B(sdata[23]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [24]) );
  MUX2_X1 \shifter_0/shift_1b_0/U79  ( .A(sdata[25]), .B(sdata[24]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [25]) );
  MUX2_X1 \shifter_0/shift_1b_0/U78  ( .A(sdata[26]), .B(sdata[25]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [26]) );
  MUX2_X1 \shifter_0/shift_1b_0/U77  ( .A(sdata[27]), .B(sdata[26]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [27]) );
  MUX2_X1 \shifter_0/shift_1b_0/U76  ( .A(sdata[28]), .B(sdata[27]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [28]) );
  MUX2_X1 \shifter_0/shift_1b_0/U75  ( .A(sdata[29]), .B(sdata[28]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [29]) );
  MUX2_X1 \shifter_0/shift_1b_0/U74  ( .A(sdata[2]), .B(sdata[1]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [2]) );
  MUX2_X1 \shifter_0/shift_1b_0/U73  ( .A(sdata[30]), .B(sdata[29]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [30]) );
  MUX2_X1 \shifter_0/shift_1b_0/U72  ( .A(sdata[31]), .B(sdata[30]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [31]) );
  MUX2_X1 \shifter_0/shift_1b_0/U71  ( .A(sdata[3]), .B(sdata[2]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [3]) );
  MUX2_X1 \shifter_0/shift_1b_0/U70  ( .A(sdata[4]), .B(sdata[3]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [4]) );
  MUX2_X1 \shifter_0/shift_1b_0/U69  ( .A(sdata[5]), .B(sdata[4]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [5]) );
  MUX2_X1 \shifter_0/shift_1b_0/U68  ( .A(sdata[6]), .B(sdata[5]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [6]) );
  MUX2_X1 \shifter_0/shift_1b_0/U67  ( .A(sdata[7]), .B(sdata[6]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [7]) );
  MUX2_X1 \shifter_0/shift_1b_0/U66  ( .A(sdata[8]), .B(sdata[7]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [8]) );
  MUX2_X1 \shifter_0/shift_1b_0/U65  ( .A(sdata[9]), .B(sdata[8]), .S(
        \shifter_0/n20 ), .Z(\shifter_0/data_1 [9]) );
  INV_X1 \shifter_0/shift_3b_0/U38  ( .A(\shifter_0/data_1 [0]), .ZN(
        \shifter_0/shift_3b_0/n38 ) );
  NOR2_X1 \shifter_0/shift_3b_0/U37  ( .A1(\shifter_0/n25 ), .A2(
        \shifter_0/shift_3b_0/n38 ), .ZN(\shifter_0/shift_3b_0/data1 [0]) );
  INV_X1 \shifter_0/shift_3b_0/U36  ( .A(\shifter_0/data_1 [1]), .ZN(
        \shifter_0/shift_3b_0/n37 ) );
  NOR2_X1 \shifter_0/shift_3b_0/U35  ( .A1(\shifter_0/n25 ), .A2(
        \shifter_0/shift_3b_0/n37 ), .ZN(\shifter_0/shift_3b_0/data1 [1]) );
  MUX2_X1 \shifter_0/shift_3b_0/U34  ( .A(\shifter_0/data_1 [5]), .B(
        \shifter_0/data_1 [3]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n10 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U33  ( .A(\shifter_0/data_1 [4]), .B(
        \shifter_0/data_1 [2]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n11 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U32  ( .A(\shifter_0/data_1 [3]), .B(
        \shifter_0/data_1 [1]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n12 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U31  ( .A(\shifter_0/data_1 [30]), .B(
        \shifter_0/data_1 [28]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n13 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U30  ( .A(\shifter_0/data_1 [2]), .B(
        \shifter_0/data_1 [0]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n14 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U29  ( .A(\shifter_0/data_1 [26]), .B(
        \shifter_0/data_1 [24]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n18 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U28  ( .A(\shifter_0/data_1 [25]), .B(
        \shifter_0/data_1 [23]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n19 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U27  ( .A(\shifter_0/data_1 [31]), .B(
        \shifter_0/data_1 [29]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n2 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U26  ( .A(\shifter_0/data_1 [24]), .B(
        \shifter_0/data_1 [22]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n20 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U25  ( .A(\shifter_0/data_1 [23]), .B(
        \shifter_0/data_1 [21]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n21 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U24  ( .A(\shifter_0/data_1 [22]), .B(
        \shifter_0/data_1 [20]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n22 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U23  ( .A(\shifter_0/data_1 [21]), .B(
        \shifter_0/data_1 [19]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n23 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U22  ( .A(\shifter_0/data_1 [20]), .B(
        \shifter_0/data_1 [18]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n24 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U21  ( .A(\shifter_0/data_1 [19]), .B(
        \shifter_0/data_1 [17]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n25 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U20  ( .A(\shifter_0/data_1 [18]), .B(
        \shifter_0/data_1 [16]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n26 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U19  ( .A(\shifter_0/data_1 [17]), .B(
        \shifter_0/data_1 [15]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n27 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U18  ( .A(\shifter_0/data_1 [16]), .B(
        \shifter_0/data_1 [14]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n28 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U17  ( .A(\shifter_0/data_1 [15]), .B(
        \shifter_0/data_1 [13]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n29 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U16  ( .A(\shifter_0/data_1 [27]), .B(
        \shifter_0/data_1 [25]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n3 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U15  ( .A(\shifter_0/data_1 [14]), .B(
        \shifter_0/data_1 [12]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n30 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U14  ( .A(\shifter_0/data_1 [13]), .B(
        \shifter_0/data_1 [11]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n31 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U13  ( .A(\shifter_0/data_1 [12]), .B(
        \shifter_0/data_1 [10]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n32 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U12  ( .A(\shifter_0/data_1 [11]), .B(
        \shifter_0/data_1 [9]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n33 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U11  ( .A(\shifter_0/data_1 [10]), .B(
        \shifter_0/data_1 [8]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n34 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U10  ( .A(\shifter_0/data_1 [28]), .B(
        \shifter_0/data_1 [26]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n4 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U9  ( .A(\shifter_0/data_1 [29]), .B(
        \shifter_0/data_1 [27]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n5 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U8  ( .A(\shifter_0/data_1 [9]), .B(
        \shifter_0/data_1 [7]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n6 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U7  ( .A(\shifter_0/data_1 [8]), .B(
        \shifter_0/data_1 [6]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n7 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U6  ( .A(\shifter_0/data_1 [7]), .B(
        \shifter_0/data_1 [5]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n8 ) );
  MUX2_X1 \shifter_0/shift_3b_0/U5  ( .A(\shifter_0/data_1 [6]), .B(
        \shifter_0/data_1 [4]), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/n9 ) );
  INV_X1 \shifter_0/shift_3b_0/U4  ( .A(1'b0), .ZN(\shifter_0/shift_3b_0/n36 )
         );
  NAND2_X1 \shifter_0/shift_3b_0/U3  ( .A1(\shifter_0/shift_3b_0/n36 ), .A2(
        \shifter_0/n4 ), .ZN(\shifter_0/shift_3b_0/n35 ) );
  MUX2_X2 \shifter_0/shift_3b_0/U2  ( .A(\shifter_0/n4 ), .B(
        \shifter_0/shift_3b_0/n35 ), .S(\shifter_0/n25 ), .Z(
        \shifter_0/shift_3b_0/shift1 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U97  ( .A(
        \shifter_0/shift_3b_0/data1 [0]), .ZN(
        \shifter_0/shift_3b_0/shift_1b_0/n33 ) );
  NOR2_X1 \shifter_0/shift_3b_0/shift_1b_0/U96  ( .A1(
        \shifter_0/shift_3b_0/shift1 ), .A2(
        \shifter_0/shift_3b_0/shift_1b_0/n33 ), .ZN(\shifter_0/data_2 [0]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U95  ( .A(
        \shifter_0/shift_3b_0/n34 ), .B(\shifter_0/shift_3b_0/n6 ), .S(
        \shifter_0/shift_3b_0/shift1 ), .Z(\shifter_0/data_2 [10]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U94  ( .A(
        \shifter_0/shift_3b_0/n33 ), .B(\shifter_0/shift_3b_0/n34 ), .S(
        \shifter_0/shift_3b_0/shift1 ), .Z(\shifter_0/data_2 [11]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U93  ( .A(
        \shifter_0/shift_3b_0/n32 ), .B(\shifter_0/shift_3b_0/n33 ), .S(
        \shifter_0/shift_3b_0/shift1 ), .Z(\shifter_0/data_2 [12]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U92  ( .A(
        \shifter_0/shift_3b_0/n31 ), .B(\shifter_0/shift_3b_0/n32 ), .S(
        \shifter_0/shift_3b_0/shift1 ), .Z(\shifter_0/data_2 [13]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U91  ( .A(
        \shifter_0/shift_3b_0/n30 ), .B(\shifter_0/shift_3b_0/n31 ), .S(
        \shifter_0/shift_3b_0/shift1 ), .Z(\shifter_0/data_2 [14]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U90  ( .A(
        \shifter_0/shift_3b_0/n29 ), .B(\shifter_0/shift_3b_0/n30 ), .S(
        \shifter_0/shift_3b_0/shift1 ), .Z(\shifter_0/data_2 [15]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U89  ( .A(
        \shifter_0/shift_3b_0/n28 ), .B(\shifter_0/shift_3b_0/n29 ), .S(
        \shifter_0/shift_3b_0/shift1 ), .Z(\shifter_0/data_2 [16]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U88  ( .A(
        \shifter_0/shift_3b_0/n27 ), .B(\shifter_0/shift_3b_0/n28 ), .S(
        \shifter_0/shift_3b_0/shift1 ), .Z(\shifter_0/data_2 [17]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U87  ( .A(
        \shifter_0/shift_3b_0/n26 ), .B(\shifter_0/shift_3b_0/n27 ), .S(
        \shifter_0/shift_3b_0/shift1 ), .Z(\shifter_0/data_2 [18]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U86  ( .A(
        \shifter_0/shift_3b_0/n25 ), .B(\shifter_0/shift_3b_0/n26 ), .S(
        \shifter_0/shift_3b_0/shift1 ), .Z(\shifter_0/data_2 [19]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U85  ( .A(
        \shifter_0/shift_3b_0/data1 [1]), .B(\shifter_0/shift_3b_0/data1 [0]), 
        .S(\shifter_0/shift_3b_0/shift1 ), .Z(\shifter_0/data_2 [1]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U84  ( .A(
        \shifter_0/shift_3b_0/n24 ), .B(\shifter_0/shift_3b_0/n25 ), .S(
        \shifter_0/shift_3b_0/shift1 ), .Z(\shifter_0/data_2 [20]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U83  ( .A(
        \shifter_0/shift_3b_0/n23 ), .B(\shifter_0/shift_3b_0/n24 ), .S(
        \shifter_0/shift_3b_0/shift1 ), .Z(\shifter_0/data_2 [21]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U82  ( .A(
        \shifter_0/shift_3b_0/n22 ), .B(\shifter_0/shift_3b_0/n23 ), .S(
        \shifter_0/shift_3b_0/shift1 ), .Z(\shifter_0/data_2 [22]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U81  ( .A(
        \shifter_0/shift_3b_0/n21 ), .B(\shifter_0/shift_3b_0/n22 ), .S(
        \shifter_0/shift_3b_0/shift1 ), .Z(\shifter_0/data_2 [23]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U80  ( .A(
        \shifter_0/shift_3b_0/n20 ), .B(\shifter_0/shift_3b_0/n21 ), .S(
        \shifter_0/shift_3b_0/shift1 ), .Z(\shifter_0/data_2 [24]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U79  ( .A(
        \shifter_0/shift_3b_0/n19 ), .B(\shifter_0/shift_3b_0/n20 ), .S(
        \shifter_0/shift_3b_0/shift1 ), .Z(\shifter_0/data_2 [25]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U78  ( .A(
        \shifter_0/shift_3b_0/n18 ), .B(\shifter_0/shift_3b_0/n19 ), .S(
        \shifter_0/shift_3b_0/shift1 ), .Z(\shifter_0/data_2 [26]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U77  ( .A(\shifter_0/shift_3b_0/n3 ), .B(\shifter_0/shift_3b_0/n18 ), .S(\shifter_0/shift_3b_0/shift1 ), .Z(
        \shifter_0/data_2 [27]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U76  ( .A(\shifter_0/shift_3b_0/n4 ), .B(\shifter_0/shift_3b_0/n3 ), .S(\shifter_0/shift_3b_0/shift1 ), .Z(
        \shifter_0/data_2 [28]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U75  ( .A(\shifter_0/shift_3b_0/n5 ), .B(\shifter_0/shift_3b_0/n4 ), .S(\shifter_0/shift_3b_0/shift1 ), .Z(
        \shifter_0/data_2 [29]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U74  ( .A(
        \shifter_0/shift_3b_0/n14 ), .B(\shifter_0/shift_3b_0/data1 [1]), .S(
        \shifter_0/shift_3b_0/shift1 ), .Z(\shifter_0/data_2 [2]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U73  ( .A(
        \shifter_0/shift_3b_0/n13 ), .B(\shifter_0/shift_3b_0/n5 ), .S(
        \shifter_0/shift_3b_0/shift1 ), .Z(\shifter_0/data_2 [30]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U72  ( .A(\shifter_0/shift_3b_0/n2 ), .B(\shifter_0/shift_3b_0/n13 ), .S(\shifter_0/shift_3b_0/shift1 ), .Z(
        \shifter_0/data_2 [31]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U71  ( .A(
        \shifter_0/shift_3b_0/n12 ), .B(\shifter_0/shift_3b_0/n14 ), .S(
        \shifter_0/shift_3b_0/shift1 ), .Z(\shifter_0/data_2 [3]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U70  ( .A(
        \shifter_0/shift_3b_0/n11 ), .B(\shifter_0/shift_3b_0/n12 ), .S(
        \shifter_0/shift_3b_0/shift1 ), .Z(\shifter_0/data_2 [4]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U69  ( .A(
        \shifter_0/shift_3b_0/n10 ), .B(\shifter_0/shift_3b_0/n11 ), .S(
        \shifter_0/shift_3b_0/shift1 ), .Z(\shifter_0/data_2 [5]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U68  ( .A(\shifter_0/shift_3b_0/n9 ), .B(\shifter_0/shift_3b_0/n10 ), .S(\shifter_0/shift_3b_0/shift1 ), .Z(
        \shifter_0/data_2 [6]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U67  ( .A(\shifter_0/shift_3b_0/n8 ), .B(\shifter_0/shift_3b_0/n9 ), .S(\shifter_0/shift_3b_0/shift1 ), .Z(
        \shifter_0/data_2 [7]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U66  ( .A(\shifter_0/shift_3b_0/n7 ), .B(\shifter_0/shift_3b_0/n8 ), .S(\shifter_0/shift_3b_0/shift1 ), .Z(
        \shifter_0/data_2 [8]) );
  MUX2_X1 \shifter_0/shift_3b_0/shift_1b_0/U65  ( .A(\shifter_0/shift_3b_0/n6 ), .B(\shifter_0/shift_3b_0/n7 ), .S(\shifter_0/shift_3b_0/shift1 ), .Z(
        \shifter_0/data_2 [9]) );
  INV_X1 \shifter_0/shift_3b_1/U38  ( .A(\shifter_0/data_2 [0]), .ZN(
        \shifter_0/shift_3b_1/n38 ) );
  NOR2_X1 \shifter_0/shift_3b_1/U37  ( .A1(\shifter_0/n24 ), .A2(
        \shifter_0/shift_3b_1/n38 ), .ZN(\shifter_0/shift_3b_1/data1 [0]) );
  INV_X1 \shifter_0/shift_3b_1/U36  ( .A(\shifter_0/data_2 [1]), .ZN(
        \shifter_0/shift_3b_1/n37 ) );
  NOR2_X1 \shifter_0/shift_3b_1/U35  ( .A1(\shifter_0/n24 ), .A2(
        \shifter_0/shift_3b_1/n37 ), .ZN(\shifter_0/shift_3b_1/data1 [1]) );
  MUX2_X1 \shifter_0/shift_3b_1/U34  ( .A(\shifter_0/data_2 [6]), .B(
        \shifter_0/data_2 [4]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n10 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U33  ( .A(\shifter_0/data_2 [5]), .B(
        \shifter_0/data_2 [3]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n11 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U32  ( .A(\shifter_0/data_2 [4]), .B(
        \shifter_0/data_2 [2]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n12 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U31  ( .A(\shifter_0/data_2 [3]), .B(
        \shifter_0/data_2 [1]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n13 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U30  ( .A(\shifter_0/data_2 [31]), .B(
        \shifter_0/data_2 [29]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n14 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U29  ( .A(\shifter_0/data_2 [2]), .B(
        \shifter_0/data_2 [0]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n16 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U28  ( .A(\shifter_0/data_2 [27]), .B(
        \shifter_0/data_2 [25]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n19 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U27  ( .A(\shifter_0/data_2 [28]), .B(
        \shifter_0/data_2 [26]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n2 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U26  ( .A(\shifter_0/data_2 [26]), .B(
        \shifter_0/data_2 [24]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n20 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U25  ( .A(\shifter_0/data_2 [25]), .B(
        \shifter_0/data_2 [23]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n21 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U24  ( .A(\shifter_0/data_2 [24]), .B(
        \shifter_0/data_2 [22]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n22 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U23  ( .A(\shifter_0/data_2 [23]), .B(
        \shifter_0/data_2 [21]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n23 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U22  ( .A(\shifter_0/data_2 [22]), .B(
        \shifter_0/data_2 [20]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n24 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U21  ( .A(\shifter_0/data_2 [21]), .B(
        \shifter_0/data_2 [19]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n25 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U20  ( .A(\shifter_0/data_2 [20]), .B(
        \shifter_0/data_2 [18]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n26 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U19  ( .A(\shifter_0/data_2 [19]), .B(
        \shifter_0/data_2 [17]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n27 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U18  ( .A(\shifter_0/data_2 [18]), .B(
        \shifter_0/data_2 [16]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n28 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U17  ( .A(\shifter_0/data_2 [17]), .B(
        \shifter_0/data_2 [15]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n29 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U16  ( .A(\shifter_0/data_2 [29]), .B(
        \shifter_0/data_2 [27]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n3 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U15  ( .A(\shifter_0/data_2 [16]), .B(
        \shifter_0/data_2 [14]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n30 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U14  ( .A(\shifter_0/data_2 [15]), .B(
        \shifter_0/data_2 [13]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n31 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U13  ( .A(\shifter_0/data_2 [14]), .B(
        \shifter_0/data_2 [12]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n32 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U12  ( .A(\shifter_0/data_2 [13]), .B(
        \shifter_0/data_2 [11]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n33 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U11  ( .A(\shifter_0/data_2 [12]), .B(
        \shifter_0/data_2 [10]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n34 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U10  ( .A(\shifter_0/data_2 [30]), .B(
        \shifter_0/data_2 [28]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n4 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U9  ( .A(\shifter_0/data_2 [11]), .B(
        \shifter_0/data_2 [9]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n5 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U8  ( .A(\shifter_0/data_2 [9]), .B(
        \shifter_0/data_2 [7]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n6 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U7  ( .A(\shifter_0/data_2 [10]), .B(
        \shifter_0/data_2 [8]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n7 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U6  ( .A(\shifter_0/data_2 [8]), .B(
        \shifter_0/data_2 [6]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n8 ) );
  MUX2_X1 \shifter_0/shift_3b_1/U5  ( .A(\shifter_0/data_2 [7]), .B(
        \shifter_0/data_2 [5]), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/n9 ) );
  INV_X1 \shifter_0/shift_3b_1/U4  ( .A(1'b0), .ZN(\shifter_0/shift_3b_1/n36 )
         );
  NAND2_X1 \shifter_0/shift_3b_1/U3  ( .A1(\shifter_0/shift_3b_1/n36 ), .A2(
        \shifter_0/n3 ), .ZN(\shifter_0/shift_3b_1/n35 ) );
  MUX2_X2 \shifter_0/shift_3b_1/U2  ( .A(\shifter_0/n3 ), .B(
        \shifter_0/shift_3b_1/n35 ), .S(\shifter_0/n24 ), .Z(
        \shifter_0/shift_3b_1/shift1 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U97  ( .A(
        \shifter_0/shift_3b_1/data1 [0]), .ZN(
        \shifter_0/shift_3b_1/shift_1b_0/n33 ) );
  NOR2_X1 \shifter_0/shift_3b_1/shift_1b_0/U96  ( .A1(
        \shifter_0/shift_3b_1/shift1 ), .A2(
        \shifter_0/shift_3b_1/shift_1b_0/n33 ), .ZN(\shifter_0/data_3 [0]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U95  ( .A(\shifter_0/shift_3b_1/n7 ), .B(\shifter_0/shift_3b_1/n6 ), .S(\shifter_0/shift_3b_1/shift1 ), .Z(
        \shifter_0/data_3 [10]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U94  ( .A(\shifter_0/shift_3b_1/n5 ), .B(\shifter_0/shift_3b_1/n7 ), .S(\shifter_0/shift_3b_1/shift1 ), .Z(
        \shifter_0/data_3 [11]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U93  ( .A(
        \shifter_0/shift_3b_1/n34 ), .B(\shifter_0/shift_3b_1/n5 ), .S(
        \shifter_0/shift_3b_1/shift1 ), .Z(\shifter_0/data_3 [12]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U92  ( .A(
        \shifter_0/shift_3b_1/n33 ), .B(\shifter_0/shift_3b_1/n34 ), .S(
        \shifter_0/shift_3b_1/shift1 ), .Z(\shifter_0/data_3 [13]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U91  ( .A(
        \shifter_0/shift_3b_1/n32 ), .B(\shifter_0/shift_3b_1/n33 ), .S(
        \shifter_0/shift_3b_1/shift1 ), .Z(\shifter_0/data_3 [14]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U90  ( .A(
        \shifter_0/shift_3b_1/n31 ), .B(\shifter_0/shift_3b_1/n32 ), .S(
        \shifter_0/shift_3b_1/shift1 ), .Z(\shifter_0/data_3 [15]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U89  ( .A(
        \shifter_0/shift_3b_1/n30 ), .B(\shifter_0/shift_3b_1/n31 ), .S(
        \shifter_0/shift_3b_1/shift1 ), .Z(\shifter_0/data_3 [16]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U88  ( .A(
        \shifter_0/shift_3b_1/n29 ), .B(\shifter_0/shift_3b_1/n30 ), .S(
        \shifter_0/shift_3b_1/shift1 ), .Z(\shifter_0/data_3 [17]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U87  ( .A(
        \shifter_0/shift_3b_1/n28 ), .B(\shifter_0/shift_3b_1/n29 ), .S(
        \shifter_0/shift_3b_1/shift1 ), .Z(\shifter_0/data_3 [18]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U86  ( .A(
        \shifter_0/shift_3b_1/n27 ), .B(\shifter_0/shift_3b_1/n28 ), .S(
        \shifter_0/shift_3b_1/shift1 ), .Z(\shifter_0/data_3 [19]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U85  ( .A(
        \shifter_0/shift_3b_1/data1 [1]), .B(\shifter_0/shift_3b_1/data1 [0]), 
        .S(\shifter_0/shift_3b_1/shift1 ), .Z(\shifter_0/data_3 [1]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U84  ( .A(
        \shifter_0/shift_3b_1/n26 ), .B(\shifter_0/shift_3b_1/n27 ), .S(
        \shifter_0/shift_3b_1/shift1 ), .Z(\shifter_0/data_3 [20]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U83  ( .A(
        \shifter_0/shift_3b_1/n25 ), .B(\shifter_0/shift_3b_1/n26 ), .S(
        \shifter_0/shift_3b_1/shift1 ), .Z(\shifter_0/data_3 [21]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U82  ( .A(
        \shifter_0/shift_3b_1/n24 ), .B(\shifter_0/shift_3b_1/n25 ), .S(
        \shifter_0/shift_3b_1/shift1 ), .Z(\shifter_0/data_3 [22]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U81  ( .A(
        \shifter_0/shift_3b_1/n23 ), .B(\shifter_0/shift_3b_1/n24 ), .S(
        \shifter_0/shift_3b_1/shift1 ), .Z(\shifter_0/data_3 [23]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U80  ( .A(
        \shifter_0/shift_3b_1/n22 ), .B(\shifter_0/shift_3b_1/n23 ), .S(
        \shifter_0/shift_3b_1/shift1 ), .Z(\shifter_0/data_3 [24]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U79  ( .A(
        \shifter_0/shift_3b_1/n21 ), .B(\shifter_0/shift_3b_1/n22 ), .S(
        \shifter_0/shift_3b_1/shift1 ), .Z(\shifter_0/data_3 [25]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U78  ( .A(
        \shifter_0/shift_3b_1/n20 ), .B(\shifter_0/shift_3b_1/n21 ), .S(
        \shifter_0/shift_3b_1/shift1 ), .Z(\shifter_0/data_3 [26]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U77  ( .A(
        \shifter_0/shift_3b_1/n19 ), .B(\shifter_0/shift_3b_1/n20 ), .S(
        \shifter_0/shift_3b_1/shift1 ), .Z(\shifter_0/data_3 [27]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U76  ( .A(\shifter_0/shift_3b_1/n2 ), .B(\shifter_0/shift_3b_1/n19 ), .S(\shifter_0/shift_3b_1/shift1 ), .Z(
        \shifter_0/data_3 [28]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U75  ( .A(\shifter_0/shift_3b_1/n3 ), .B(\shifter_0/shift_3b_1/n2 ), .S(\shifter_0/shift_3b_1/shift1 ), .Z(
        \shifter_0/data_3 [29]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U74  ( .A(
        \shifter_0/shift_3b_1/n16 ), .B(\shifter_0/shift_3b_1/data1 [1]), .S(
        \shifter_0/shift_3b_1/shift1 ), .Z(\shifter_0/data_3 [2]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U73  ( .A(\shifter_0/shift_3b_1/n4 ), .B(\shifter_0/shift_3b_1/n3 ), .S(\shifter_0/shift_3b_1/shift1 ), .Z(
        \shifter_0/data_3 [30]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U72  ( .A(
        \shifter_0/shift_3b_1/n14 ), .B(\shifter_0/shift_3b_1/n4 ), .S(
        \shifter_0/shift_3b_1/shift1 ), .Z(\shifter_0/data_3 [31]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U71  ( .A(
        \shifter_0/shift_3b_1/n13 ), .B(\shifter_0/shift_3b_1/n16 ), .S(
        \shifter_0/shift_3b_1/shift1 ), .Z(\shifter_0/data_3 [3]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U70  ( .A(
        \shifter_0/shift_3b_1/n12 ), .B(\shifter_0/shift_3b_1/n13 ), .S(
        \shifter_0/shift_3b_1/shift1 ), .Z(\shifter_0/data_3 [4]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U69  ( .A(
        \shifter_0/shift_3b_1/n11 ), .B(\shifter_0/shift_3b_1/n12 ), .S(
        \shifter_0/shift_3b_1/shift1 ), .Z(\shifter_0/data_3 [5]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U68  ( .A(
        \shifter_0/shift_3b_1/n10 ), .B(\shifter_0/shift_3b_1/n11 ), .S(
        \shifter_0/shift_3b_1/shift1 ), .Z(\shifter_0/data_3 [6]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U67  ( .A(\shifter_0/shift_3b_1/n9 ), .B(\shifter_0/shift_3b_1/n10 ), .S(\shifter_0/shift_3b_1/shift1 ), .Z(
        \shifter_0/data_3 [7]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U66  ( .A(\shifter_0/shift_3b_1/n8 ), .B(\shifter_0/shift_3b_1/n9 ), .S(\shifter_0/shift_3b_1/shift1 ), .Z(
        \shifter_0/data_3 [8]) );
  MUX2_X1 \shifter_0/shift_3b_1/shift_1b_0/U65  ( .A(\shifter_0/shift_3b_1/n6 ), .B(\shifter_0/shift_3b_1/n8 ), .S(\shifter_0/shift_3b_1/shift1 ), .Z(
        \shifter_0/data_3 [9]) );
  INV_X1 \shifter_0/shift_7b_0/U46  ( .A(\shifter_0/data_3 [0]), .ZN(
        \shifter_0/shift_7b_0/n48 ) );
  NOR2_X1 \shifter_0/shift_7b_0/U45  ( .A1(\shifter_0/n21 ), .A2(
        \shifter_0/shift_7b_0/n48 ), .ZN(\shifter_0/shift_7b_0/data1 [0]) );
  INV_X1 \shifter_0/shift_7b_0/U44  ( .A(\shifter_0/data_3 [1]), .ZN(
        \shifter_0/shift_7b_0/n47 ) );
  NOR2_X1 \shifter_0/shift_7b_0/U43  ( .A1(\shifter_0/n21 ), .A2(
        \shifter_0/shift_7b_0/n47 ), .ZN(\shifter_0/shift_7b_0/data1 [1]) );
  INV_X1 \shifter_0/shift_7b_0/U42  ( .A(\shifter_0/data_3 [2]), .ZN(
        \shifter_0/shift_7b_0/n46 ) );
  NOR2_X1 \shifter_0/shift_7b_0/U41  ( .A1(\shifter_0/n21 ), .A2(
        \shifter_0/shift_7b_0/n46 ), .ZN(\shifter_0/shift_7b_0/data1 [2]) );
  INV_X1 \shifter_0/shift_7b_0/U40  ( .A(\shifter_0/data_3 [3]), .ZN(
        \shifter_0/shift_7b_0/n45 ) );
  NOR2_X1 \shifter_0/shift_7b_0/U39  ( .A1(\shifter_0/n21 ), .A2(
        \shifter_0/shift_7b_0/n45 ), .ZN(\shifter_0/shift_7b_0/data1 [3]) );
  MUX2_X1 \shifter_0/shift_7b_0/U38  ( .A(\shifter_0/data_3 [30]), .B(
        \shifter_0/data_3 [26]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n10 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U37  ( .A(\shifter_0/data_3 [13]), .B(
        \shifter_0/data_3 [9]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n11 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U36  ( .A(\shifter_0/data_3 [9]), .B(
        \shifter_0/data_3 [5]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n12 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U35  ( .A(\shifter_0/data_3 [12]), .B(
        \shifter_0/data_3 [8]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n13 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U34  ( .A(\shifter_0/data_3 [8]), .B(
        \shifter_0/data_3 [4]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n14 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U33  ( .A(\shifter_0/data_3 [11]), .B(
        \shifter_0/data_3 [7]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n15 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U32  ( .A(\shifter_0/data_3 [7]), .B(
        \shifter_0/data_3 [3]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n16 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U31  ( .A(\shifter_0/data_3 [10]), .B(
        \shifter_0/data_3 [6]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n17 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U30  ( .A(\shifter_0/data_3 [6]), .B(
        \shifter_0/data_3 [2]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n18 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U29  ( .A(\shifter_0/data_3 [5]), .B(
        \shifter_0/data_3 [1]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n19 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U28  ( .A(\shifter_0/data_3 [4]), .B(
        \shifter_0/data_3 [0]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n20 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U27  ( .A(\shifter_0/data_3 [31]), .B(
        \shifter_0/data_3 [27]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n21 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U26  ( .A(\shifter_0/data_3 [23]), .B(
        \shifter_0/data_3 [19]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n29 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U25  ( .A(\shifter_0/data_3 [22]), .B(
        \shifter_0/data_3 [18]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n30 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U24  ( .A(\shifter_0/data_3 [21]), .B(
        \shifter_0/data_3 [17]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n31 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U23  ( .A(\shifter_0/data_3 [20]), .B(
        \shifter_0/data_3 [16]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n32 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U22  ( .A(\shifter_0/data_3 [19]), .B(
        \shifter_0/data_3 [15]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n33 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U21  ( .A(\shifter_0/data_3 [18]), .B(
        \shifter_0/data_3 [14]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n34 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U20  ( .A(\shifter_0/data_3 [17]), .B(
        \shifter_0/data_3 [13]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n35 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U19  ( .A(\shifter_0/data_3 [16]), .B(
        \shifter_0/data_3 [12]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n36 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U18  ( .A(\shifter_0/data_3 [15]), .B(
        \shifter_0/data_3 [11]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n37 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U17  ( .A(\shifter_0/data_3 [14]), .B(
        \shifter_0/data_3 [10]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n38 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U16  ( .A(\shifter_0/data_3 [24]), .B(
        \shifter_0/data_3 [20]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n4 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U15  ( .A(\shifter_0/data_3 [25]), .B(
        \shifter_0/data_3 [21]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n5 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U14  ( .A(\shifter_0/data_3 [26]), .B(
        \shifter_0/data_3 [22]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n6 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U13  ( .A(\shifter_0/data_3 [27]), .B(
        \shifter_0/data_3 [23]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n7 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U12  ( .A(\shifter_0/data_3 [28]), .B(
        \shifter_0/data_3 [24]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n8 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U11  ( .A(\shifter_0/data_3 [29]), .B(
        \shifter_0/data_3 [25]), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/n9 ) );
  INV_X1 \shifter_0/shift_7b_0/U10  ( .A(1'b0), .ZN(\shifter_0/shift_7b_0/n44 ) );
  NAND2_X1 \shifter_0/shift_7b_0/U9  ( .A1(\shifter_0/shift_7b_0/n44 ), .A2(
        shifted_o[3]), .ZN(\shifter_0/shift_7b_0/n43 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U8  ( .A(shifted_o[3]), .B(
        \shifter_0/shift_7b_0/n43 ), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/shift1 [0]) );
  INV_X1 \shifter_0/shift_7b_0/U7  ( .A(1'b0), .ZN(\shifter_0/shift_7b_0/n42 )
         );
  NAND2_X1 \shifter_0/shift_7b_0/U6  ( .A1(\shifter_0/shift_7b_0/n42 ), .A2(
        \shifter_0/n1 ), .ZN(\shifter_0/shift_7b_0/n41 ) );
  INV_X1 \shifter_0/shift_7b_0/U5  ( .A(1'b0), .ZN(\shifter_0/shift_7b_0/n40 )
         );
  NAND2_X1 \shifter_0/shift_7b_0/U4  ( .A1(\shifter_0/shift_7b_0/n40 ), .A2(
        \shifter_0/n2 ), .ZN(\shifter_0/shift_7b_0/n39 ) );
  MUX2_X1 \shifter_0/shift_7b_0/U3  ( .A(\shifter_0/n2 ), .B(
        \shifter_0/shift_7b_0/n39 ), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/shift1 [2]) );
  MUX2_X2 \shifter_0/shift_7b_0/U2  ( .A(\shifter_0/n1 ), .B(
        \shifter_0/shift_7b_0/n41 ), .S(\shifter_0/n21 ), .Z(
        \shifter_0/shift_7b_0/shift1 [1]) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U38  ( .A(
        \shifter_0/shift_7b_0/data1 [0]), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n38 ) );
  NOR2_X1 \shifter_0/shift_7b_0/shift_3b_0/U37  ( .A1(
        \shifter_0/shift_7b_0/shift1 [1]), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n38 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/data1 [0]) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U36  ( .A(
        \shifter_0/shift_7b_0/data1 [1]), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ) );
  NOR2_X1 \shifter_0/shift_7b_0/shift_3b_0/U35  ( .A1(
        \shifter_0/shift_7b_0/shift1 [1]), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/data1 [1]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U34  ( .A(
        \shifter_0/shift_7b_0/n38 ), .B(\shifter_0/shift_7b_0/n13 ), .S(
        \shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n10 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U33  ( .A(
        \shifter_0/shift_7b_0/n17 ), .B(\shifter_0/shift_7b_0/n14 ), .S(
        \shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n11 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U32  ( .A(
        \shifter_0/shift_7b_0/n14 ), .B(\shifter_0/shift_7b_0/n18 ), .S(
        \shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n12 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U31  ( .A(
        \shifter_0/shift_7b_0/n16 ), .B(\shifter_0/shift_7b_0/n19 ), .S(
        \shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n13 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U30  ( .A(
        \shifter_0/shift_7b_0/n18 ), .B(\shifter_0/shift_7b_0/n20 ), .S(
        \shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n14 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U29  ( .A(
        \shifter_0/shift_7b_0/n19 ), .B(\shifter_0/shift_7b_0/data1 [3]), .S(
        \shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n15 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U28  ( .A(
        \shifter_0/shift_7b_0/n20 ), .B(\shifter_0/shift_7b_0/data1 [2]), .S(
        \shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n16 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U27  ( .A(
        \shifter_0/shift_7b_0/data1 [3]), .B(\shifter_0/shift_7b_0/data1 [1]), 
        .S(\shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n17 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U26  ( .A(
        \shifter_0/shift_7b_0/n21 ), .B(\shifter_0/shift_7b_0/n9 ), .S(
        \shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n18 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U25  ( .A(\shifter_0/shift_7b_0/n8 ), .B(\shifter_0/shift_7b_0/n6 ), .S(\shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n2 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U24  ( .A(
        \shifter_0/shift_7b_0/data1 [2]), .B(\shifter_0/shift_7b_0/data1 [0]), 
        .S(\shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n20 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U23  ( .A(\shifter_0/shift_7b_0/n7 ), .B(\shifter_0/shift_7b_0/n5 ), .S(\shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n23 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U22  ( .A(\shifter_0/shift_7b_0/n6 ), .B(\shifter_0/shift_7b_0/n4 ), .S(\shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n24 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U21  ( .A(\shifter_0/shift_7b_0/n5 ), .B(\shifter_0/shift_7b_0/n29 ), .S(\shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n25 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U20  ( .A(\shifter_0/shift_7b_0/n4 ), .B(\shifter_0/shift_7b_0/n30 ), .S(\shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n26 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U19  ( .A(
        \shifter_0/shift_7b_0/n29 ), .B(\shifter_0/shift_7b_0/n31 ), .S(
        \shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n27 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U18  ( .A(
        \shifter_0/shift_7b_0/n30 ), .B(\shifter_0/shift_7b_0/n32 ), .S(
        \shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n28 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U17  ( .A(
        \shifter_0/shift_7b_0/n31 ), .B(\shifter_0/shift_7b_0/n33 ), .S(
        \shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n29 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U16  ( .A(\shifter_0/shift_7b_0/n9 ), .B(\shifter_0/shift_7b_0/n7 ), .S(\shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n3 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U15  ( .A(
        \shifter_0/shift_7b_0/n32 ), .B(\shifter_0/shift_7b_0/n34 ), .S(
        \shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n30 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U14  ( .A(
        \shifter_0/shift_7b_0/n33 ), .B(\shifter_0/shift_7b_0/n35 ), .S(
        \shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n31 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U13  ( .A(
        \shifter_0/shift_7b_0/n34 ), .B(\shifter_0/shift_7b_0/n36 ), .S(
        \shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n32 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U12  ( .A(
        \shifter_0/shift_7b_0/n35 ), .B(\shifter_0/shift_7b_0/n37 ), .S(
        \shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n33 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U11  ( .A(
        \shifter_0/shift_7b_0/n36 ), .B(\shifter_0/shift_7b_0/n38 ), .S(
        \shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n34 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U10  ( .A(
        \shifter_0/shift_7b_0/n10 ), .B(\shifter_0/shift_7b_0/n8 ), .S(
        \shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n4 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U9  ( .A(\shifter_0/shift_7b_0/n11 ), .B(\shifter_0/shift_7b_0/n15 ), .S(\shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n5 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U8  ( .A(\shifter_0/shift_7b_0/n37 ), .B(\shifter_0/shift_7b_0/n11 ), .S(\shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n6 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U7  ( .A(\shifter_0/shift_7b_0/n15 ), .B(\shifter_0/shift_7b_0/n12 ), .S(\shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n7 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U6  ( .A(\shifter_0/shift_7b_0/n12 ), .B(\shifter_0/shift_7b_0/n16 ), .S(\shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n8 ) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/U5  ( .A(\shifter_0/shift_7b_0/n13 ), .B(\shifter_0/shift_7b_0/n17 ), .S(\shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n9 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U4  ( .A(
        \shifter_0/shift_7b_0/shift1 [0]), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n36 ) );
  NAND2_X1 \shifter_0/shift_7b_0/shift_3b_0/U3  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_7b_0/shift1 [2]), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n35 ) );
  MUX2_X2 \shifter_0/shift_7b_0/shift_3b_0/U2  ( .A(
        \shifter_0/shift_7b_0/shift1 [2]), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n35 ), .S(
        \shifter_0/shift_7b_0/shift1 [1]), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U97  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/data1 [0]), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n33 ) );
  NOR2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U96  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n33 ), .ZN(sdata_o[0]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U95  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n11 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n8 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[10]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U94  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n7 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n11 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[11]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U93  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n9 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n7 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[12]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U92  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n5 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n9 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[13]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U91  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n10 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n5 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[14]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U90  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n6 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n10 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[15]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U89  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n34 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n6 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[16]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U88  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n33 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n34 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[17]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U87  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n32 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n33 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[18]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U86  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n31 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n32 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[19]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U85  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/data1 [1]), .B(
        \shifter_0/shift_7b_0/shift_3b_0/data1 [0]), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[1]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U84  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n30 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n31 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[20]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U83  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n29 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n30 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[21]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U82  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n28 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n29 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[22]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U81  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n27 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n28 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[23]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U80  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n26 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n27 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[24]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U79  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n25 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n26 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[25]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U78  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n24 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n25 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[26]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U77  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n23 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n24 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[27]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U76  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n2 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n23 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[28]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U75  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n3 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n2 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[29]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U74  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n20 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/data1 [1]), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[2]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U73  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n4 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n3 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[30]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U72  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n18 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n4 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[31]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U71  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n17 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n20 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[3]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U70  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n16 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n17 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[4]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U69  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n15 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n16 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[5]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U68  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n14 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n15 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[6]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U67  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n13 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n14 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[7]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U66  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n12 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n13 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[8]) );
  MUX2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U65  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n8 ), .B(
        \shifter_0/shift_7b_0/shift_3b_0/n12 ), .S(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(sdata_o[9]) );
  XOR2_X1 \adder_0/U32  ( .A(reg_carry), .B(\adder_0/P0[0] ), .Z(sum[0]) );
  XOR2_X1 \adder_0/U31  ( .A(\adder_0/P0[10] ), .B(\adder_0/G6_9 ), .Z(sum[10]) );
  XOR2_X1 \adder_0/U30  ( .A(\adder_0/P0[11] ), .B(\adder_0/G4[5] ), .Z(
        sum[11]) );
  XOR2_X1 \adder_0/U29  ( .A(\adder_0/P0[12] ), .B(\adder_0/G6_11 ), .Z(
        sum[12]) );
  XOR2_X1 \adder_0/U28  ( .A(\adder_0/P0[13] ), .B(\adder_0/G4[6] ), .Z(
        sum[13]) );
  XOR2_X1 \adder_0/U27  ( .A(\adder_0/P0[14] ), .B(\adder_0/G6_13 ), .Z(
        sum[14]) );
  XOR2_X1 \adder_0/U26  ( .A(\adder_0/P0[15] ), .B(\adder_0/G4[7] ), .Z(
        sum[15]) );
  XOR2_X1 \adder_0/U25  ( .A(\adder_0/P0[16] ), .B(\adder_0/G6_15 ), .Z(
        sum[16]) );
  XOR2_X1 \adder_0/U24  ( .A(\adder_0/P0[17] ), .B(\adder_0/G5[8] ), .Z(
        sum[17]) );
  XOR2_X1 \adder_0/U23  ( .A(\adder_0/P0[18] ), .B(\adder_0/G6_17 ), .Z(
        sum[18]) );
  XOR2_X1 \adder_0/U22  ( .A(\adder_0/P0[19] ), .B(\adder_0/G5[9] ), .Z(
        sum[19]) );
  XOR2_X1 \adder_0/U21  ( .A(\adder_0/P0[1] ), .B(\adder_0/G1[0] ), .Z(sum[1])
         );
  XOR2_X1 \adder_0/U20  ( .A(\adder_0/P0[20] ), .B(\adder_0/G6_19 ), .Z(
        sum[20]) );
  XOR2_X1 \adder_0/U19  ( .A(\adder_0/P0[21] ), .B(\adder_0/G5[10] ), .Z(
        sum[21]) );
  XOR2_X1 \adder_0/U18  ( .A(\adder_0/P0[22] ), .B(\adder_0/G6_21 ), .Z(
        sum[22]) );
  XOR2_X1 \adder_0/U17  ( .A(\adder_0/P0[23] ), .B(\adder_0/G5[11] ), .Z(
        sum[23]) );
  XOR2_X1 \adder_0/U16  ( .A(\adder_0/P0[24] ), .B(\adder_0/G6_23 ), .Z(
        sum[24]) );
  XOR2_X1 \adder_0/U15  ( .A(\adder_0/P0[25] ), .B(\adder_0/G5[12] ), .Z(
        sum[25]) );
  XOR2_X1 \adder_0/U14  ( .A(\adder_0/P0[26] ), .B(\adder_0/G6_25 ), .Z(
        sum[26]) );
  XOR2_X1 \adder_0/U13  ( .A(\adder_0/P0[27] ), .B(\adder_0/G5[13] ), .Z(
        sum[27]) );
  XOR2_X1 \adder_0/U12  ( .A(\adder_0/P0[28] ), .B(\adder_0/G6_27 ), .Z(
        sum[28]) );
  XOR2_X1 \adder_0/U11  ( .A(\adder_0/P0[29] ), .B(\adder_0/G5[14] ), .Z(
        sum[29]) );
  XOR2_X1 \adder_0/U10  ( .A(\adder_0/P0[2] ), .B(\adder_0/G6_1 ), .Z(sum[2])
         );
  XOR2_X1 \adder_0/U9  ( .A(\adder_0/P0[30] ), .B(\adder_0/G6_29_ ), .Z(
        sum[30]) );
  XOR2_X1 \adder_0/U8  ( .A(\adder_0/P0[31] ), .B(\adder_0/G5[15] ), .Z(
        sum[31]) );
  XOR2_X1 \adder_0/U7  ( .A(\adder_0/P0[3] ), .B(\adder_0/G2[1] ), .Z(sum[3])
         );
  XOR2_X1 \adder_0/U6  ( .A(\adder_0/P0[4] ), .B(\adder_0/G6_3 ), .Z(sum[4])
         );
  XOR2_X1 \adder_0/U5  ( .A(\adder_0/P0[5] ), .B(\adder_0/G3[2] ), .Z(sum[5])
         );
  XOR2_X1 \adder_0/U4  ( .A(\adder_0/P0[6] ), .B(\adder_0/G6_5 ), .Z(sum[6])
         );
  XOR2_X1 \adder_0/U3  ( .A(\adder_0/P0[7] ), .B(\adder_0/G3[3] ), .Z(sum[7])
         );
  XOR2_X1 \adder_0/U2  ( .A(\adder_0/P0[8] ), .B(\adder_0/G6_7 ), .Z(sum[8])
         );
  XOR2_X1 \adder_0/U1  ( .A(\adder_0/P0[9] ), .B(\adder_0/G4[4] ), .Z(sum[9])
         );
  AND2_X1 \adder_0/operator_A_0/U2  ( .A1(reg_b[0]), .A2(reg_a[0]), .ZN(
        \adder_0/G0[0] ) );
  XOR2_X1 \adder_0/operator_A_0/U1  ( .A(reg_b[0]), .B(reg_a[0]), .Z(
        \adder_0/P0[0] ) );
  AND2_X1 \adder_0/operator_A_1/U2  ( .A1(reg_b[1]), .A2(reg_a[1]), .ZN(
        \adder_0/G0[1] ) );
  XOR2_X1 \adder_0/operator_A_1/U1  ( .A(reg_b[1]), .B(reg_a[1]), .Z(
        \adder_0/P0[1] ) );
  AND2_X1 \adder_0/operator_A_2/U2  ( .A1(reg_b[2]), .A2(reg_a[2]), .ZN(
        \adder_0/G0[2] ) );
  XOR2_X1 \adder_0/operator_A_2/U1  ( .A(reg_b[2]), .B(reg_a[2]), .Z(
        \adder_0/P0[2] ) );
  AND2_X1 \adder_0/operator_A_3/U2  ( .A1(reg_b[3]), .A2(reg_a[3]), .ZN(
        \adder_0/G0[3] ) );
  XOR2_X1 \adder_0/operator_A_3/U1  ( .A(reg_b[3]), .B(reg_a[3]), .Z(
        \adder_0/P0[3] ) );
  AND2_X1 \adder_0/operator_A_4/U2  ( .A1(reg_b[4]), .A2(reg_a[4]), .ZN(
        \adder_0/G0[4] ) );
  XOR2_X1 \adder_0/operator_A_4/U1  ( .A(reg_b[4]), .B(reg_a[4]), .Z(
        \adder_0/P0[4] ) );
  AND2_X1 \adder_0/operator_A_5/U2  ( .A1(reg_b[5]), .A2(reg_a[5]), .ZN(
        \adder_0/G0[5] ) );
  XOR2_X1 \adder_0/operator_A_5/U1  ( .A(reg_b[5]), .B(reg_a[5]), .Z(
        \adder_0/P0[5] ) );
  AND2_X1 \adder_0/operator_A_6/U2  ( .A1(reg_b[6]), .A2(reg_a[6]), .ZN(
        \adder_0/G0[6] ) );
  XOR2_X1 \adder_0/operator_A_6/U1  ( .A(reg_b[6]), .B(reg_a[6]), .Z(
        \adder_0/P0[6] ) );
  AND2_X1 \adder_0/operator_A_7/U2  ( .A1(reg_b[7]), .A2(reg_a[7]), .ZN(
        \adder_0/G0[7] ) );
  XOR2_X1 \adder_0/operator_A_7/U1  ( .A(reg_b[7]), .B(reg_a[7]), .Z(
        \adder_0/P0[7] ) );
  AND2_X1 \adder_0/operator_A_8/U2  ( .A1(reg_b[8]), .A2(reg_a[8]), .ZN(
        \adder_0/G0[8] ) );
  XOR2_X1 \adder_0/operator_A_8/U1  ( .A(reg_b[8]), .B(reg_a[8]), .Z(
        \adder_0/P0[8] ) );
  AND2_X1 \adder_0/operator_A_9/U2  ( .A1(reg_b[9]), .A2(reg_a[9]), .ZN(
        \adder_0/G0[9] ) );
  XOR2_X1 \adder_0/operator_A_9/U1  ( .A(reg_b[9]), .B(reg_a[9]), .Z(
        \adder_0/P0[9] ) );
  AND2_X1 \adder_0/operator_A_10/U2  ( .A1(reg_b[10]), .A2(reg_a[10]), .ZN(
        \adder_0/G0[10] ) );
  XOR2_X1 \adder_0/operator_A_10/U1  ( .A(reg_b[10]), .B(reg_a[10]), .Z(
        \adder_0/P0[10] ) );
  AND2_X1 \adder_0/operator_A_11/U2  ( .A1(reg_b[11]), .A2(reg_a[11]), .ZN(
        \adder_0/G0[11] ) );
  XOR2_X1 \adder_0/operator_A_11/U1  ( .A(reg_b[11]), .B(reg_a[11]), .Z(
        \adder_0/P0[11] ) );
  AND2_X1 \adder_0/operator_A_12/U2  ( .A1(reg_b[12]), .A2(reg_a[12]), .ZN(
        \adder_0/G0[12] ) );
  XOR2_X1 \adder_0/operator_A_12/U1  ( .A(reg_b[12]), .B(reg_a[12]), .Z(
        \adder_0/P0[12] ) );
  AND2_X1 \adder_0/operator_A_13/U2  ( .A1(reg_b[13]), .A2(reg_a[13]), .ZN(
        \adder_0/G0[13] ) );
  XOR2_X1 \adder_0/operator_A_13/U1  ( .A(reg_b[13]), .B(reg_a[13]), .Z(
        \adder_0/P0[13] ) );
  AND2_X1 \adder_0/operator_A_14/U2  ( .A1(reg_b[14]), .A2(reg_a[14]), .ZN(
        \adder_0/G0[14] ) );
  XOR2_X1 \adder_0/operator_A_14/U1  ( .A(reg_b[14]), .B(reg_a[14]), .Z(
        \adder_0/P0[14] ) );
  AND2_X1 \adder_0/operator_A_15/U2  ( .A1(reg_b[15]), .A2(reg_a[15]), .ZN(
        \adder_0/G0[15] ) );
  XOR2_X1 \adder_0/operator_A_15/U1  ( .A(reg_b[15]), .B(reg_a[15]), .Z(
        \adder_0/P0[15] ) );
  AND2_X1 \adder_0/operator_A_16/U2  ( .A1(reg_b[16]), .A2(reg_a[16]), .ZN(
        \adder_0/G0[16] ) );
  XOR2_X1 \adder_0/operator_A_16/U1  ( .A(reg_b[16]), .B(reg_a[16]), .Z(
        \adder_0/P0[16] ) );
  AND2_X1 \adder_0/operator_A_17/U2  ( .A1(reg_b[17]), .A2(reg_a[17]), .ZN(
        \adder_0/G0[17] ) );
  XOR2_X1 \adder_0/operator_A_17/U1  ( .A(reg_b[17]), .B(reg_a[17]), .Z(
        \adder_0/P0[17] ) );
  AND2_X1 \adder_0/operator_A_18/U2  ( .A1(reg_b[18]), .A2(reg_a[18]), .ZN(
        \adder_0/G0[18] ) );
  XOR2_X1 \adder_0/operator_A_18/U1  ( .A(reg_b[18]), .B(reg_a[18]), .Z(
        \adder_0/P0[18] ) );
  AND2_X1 \adder_0/operator_A_19/U2  ( .A1(reg_b[19]), .A2(reg_a[19]), .ZN(
        \adder_0/G0[19] ) );
  XOR2_X1 \adder_0/operator_A_19/U1  ( .A(reg_b[19]), .B(reg_a[19]), .Z(
        \adder_0/P0[19] ) );
  AND2_X1 \adder_0/operator_A_20/U2  ( .A1(reg_b[20]), .A2(reg_a[20]), .ZN(
        \adder_0/G0[20] ) );
  XOR2_X1 \adder_0/operator_A_20/U1  ( .A(reg_b[20]), .B(reg_a[20]), .Z(
        \adder_0/P0[20] ) );
  AND2_X1 \adder_0/operator_A_21/U2  ( .A1(reg_b[21]), .A2(reg_a[21]), .ZN(
        \adder_0/G0[21] ) );
  XOR2_X1 \adder_0/operator_A_21/U1  ( .A(reg_b[21]), .B(reg_a[21]), .Z(
        \adder_0/P0[21] ) );
  AND2_X1 \adder_0/operator_A_22/U2  ( .A1(reg_b[22]), .A2(reg_a[22]), .ZN(
        \adder_0/G0[22] ) );
  XOR2_X1 \adder_0/operator_A_22/U1  ( .A(reg_b[22]), .B(reg_a[22]), .Z(
        \adder_0/P0[22] ) );
  AND2_X1 \adder_0/operator_A_23/U2  ( .A1(reg_b[23]), .A2(reg_a[23]), .ZN(
        \adder_0/G0[23] ) );
  XOR2_X1 \adder_0/operator_A_23/U1  ( .A(reg_b[23]), .B(reg_a[23]), .Z(
        \adder_0/P0[23] ) );
  AND2_X1 \adder_0/operator_A_24/U2  ( .A1(reg_b[24]), .A2(reg_a[24]), .ZN(
        \adder_0/G0[24] ) );
  XOR2_X1 \adder_0/operator_A_24/U1  ( .A(reg_b[24]), .B(reg_a[24]), .Z(
        \adder_0/P0[24] ) );
  AND2_X1 \adder_0/operator_A_25/U2  ( .A1(reg_b[25]), .A2(reg_a[25]), .ZN(
        \adder_0/G0[25] ) );
  XOR2_X1 \adder_0/operator_A_25/U1  ( .A(reg_b[25]), .B(reg_a[25]), .Z(
        \adder_0/P0[25] ) );
  AND2_X1 \adder_0/operator_A_26/U2  ( .A1(reg_b[26]), .A2(reg_a[26]), .ZN(
        \adder_0/G0[26] ) );
  XOR2_X1 \adder_0/operator_A_26/U1  ( .A(reg_b[26]), .B(reg_a[26]), .Z(
        \adder_0/P0[26] ) );
  AND2_X1 \adder_0/operator_A_27/U2  ( .A1(reg_b[27]), .A2(reg_a[27]), .ZN(
        \adder_0/G0[27] ) );
  XOR2_X1 \adder_0/operator_A_27/U1  ( .A(reg_b[27]), .B(reg_a[27]), .Z(
        \adder_0/P0[27] ) );
  AND2_X1 \adder_0/operator_A_28/U2  ( .A1(reg_b[28]), .A2(reg_a[28]), .ZN(
        \adder_0/G0[28] ) );
  XOR2_X1 \adder_0/operator_A_28/U1  ( .A(reg_b[28]), .B(reg_a[28]), .Z(
        \adder_0/P0[28] ) );
  AND2_X1 \adder_0/operator_A_29/U2  ( .A1(reg_b[29]), .A2(reg_a[29]), .ZN(
        \adder_0/G0[29] ) );
  XOR2_X1 \adder_0/operator_A_29/U1  ( .A(reg_b[29]), .B(reg_a[29]), .Z(
        \adder_0/P0[29] ) );
  AND2_X1 \adder_0/operator_A_30/U2  ( .A1(reg_b[30]), .A2(reg_a[30]), .ZN(
        \adder_0/G0[30] ) );
  XOR2_X1 \adder_0/operator_A_30/U1  ( .A(reg_b[30]), .B(reg_a[30]), .Z(
        \adder_0/P0[30] ) );
  AND2_X1 \adder_0/operator_A_31/U2  ( .A1(reg_b[31]), .A2(reg_a[31]), .ZN(
        \adder_0/G0[31] ) );
  XOR2_X1 \adder_0/operator_A_31/U1  ( .A(reg_b[31]), .B(reg_a[31]), .Z(
        \adder_0/P0[31] ) );
  AOI21_X1 \adder_0/operator_C_stage_1_0/U2  ( .B1(\adder_0/P0[0] ), .B2(
        reg_carry), .A(\adder_0/G0[0] ), .ZN(\adder_0/operator_C_stage_1_0/n3 ) );
  INV_X1 \adder_0/operator_C_stage_1_0/U1  ( .A(
        \adder_0/operator_C_stage_1_0/n3 ), .ZN(\adder_0/G1[0] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_1/U3  ( .B1(\adder_0/G0[1] ), .B2(
        \adder_0/P0[2] ), .A(\adder_0/G0[2] ), .ZN(
        \adder_0/operator_B_stage_1_1/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_1/U2  ( .A(
        \adder_0/operator_B_stage_1_1/n3 ), .ZN(\adder_0/G1[1] ) );
  AND2_X1 \adder_0/operator_B_stage_1_1/U1  ( .A1(\adder_0/P0[1] ), .A2(
        \adder_0/P0[2] ), .ZN(\adder_0/P1[1] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_2/U3  ( .B1(\adder_0/G0[3] ), .B2(
        \adder_0/P0[4] ), .A(\adder_0/G0[4] ), .ZN(
        \adder_0/operator_B_stage_1_2/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_2/U2  ( .A(
        \adder_0/operator_B_stage_1_2/n3 ), .ZN(\adder_0/G1[2] ) );
  AND2_X1 \adder_0/operator_B_stage_1_2/U1  ( .A1(\adder_0/P0[3] ), .A2(
        \adder_0/P0[4] ), .ZN(\adder_0/P1[2] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_3/U3  ( .B1(\adder_0/G0[5] ), .B2(
        \adder_0/P0[6] ), .A(\adder_0/G0[6] ), .ZN(
        \adder_0/operator_B_stage_1_3/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_3/U2  ( .A(
        \adder_0/operator_B_stage_1_3/n3 ), .ZN(\adder_0/G1[3] ) );
  AND2_X1 \adder_0/operator_B_stage_1_3/U1  ( .A1(\adder_0/P0[5] ), .A2(
        \adder_0/P0[6] ), .ZN(\adder_0/P1[3] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_4/U3  ( .B1(\adder_0/G0[7] ), .B2(
        \adder_0/P0[8] ), .A(\adder_0/G0[8] ), .ZN(
        \adder_0/operator_B_stage_1_4/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_4/U2  ( .A(
        \adder_0/operator_B_stage_1_4/n3 ), .ZN(\adder_0/G1[4] ) );
  AND2_X1 \adder_0/operator_B_stage_1_4/U1  ( .A1(\adder_0/P0[7] ), .A2(
        \adder_0/P0[8] ), .ZN(\adder_0/P1[4] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_5/U3  ( .B1(\adder_0/G0[9] ), .B2(
        \adder_0/P0[10] ), .A(\adder_0/G0[10] ), .ZN(
        \adder_0/operator_B_stage_1_5/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_5/U2  ( .A(
        \adder_0/operator_B_stage_1_5/n3 ), .ZN(\adder_0/G1[5] ) );
  AND2_X1 \adder_0/operator_B_stage_1_5/U1  ( .A1(\adder_0/P0[9] ), .A2(
        \adder_0/P0[10] ), .ZN(\adder_0/P1[5] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_6/U3  ( .B1(\adder_0/G0[11] ), .B2(
        \adder_0/P0[12] ), .A(\adder_0/G0[12] ), .ZN(
        \adder_0/operator_B_stage_1_6/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_6/U2  ( .A(
        \adder_0/operator_B_stage_1_6/n3 ), .ZN(\adder_0/G1[6] ) );
  AND2_X1 \adder_0/operator_B_stage_1_6/U1  ( .A1(\adder_0/P0[11] ), .A2(
        \adder_0/P0[12] ), .ZN(\adder_0/P1[6] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_7/U3  ( .B1(\adder_0/G0[13] ), .B2(
        \adder_0/P0[14] ), .A(\adder_0/G0[14] ), .ZN(
        \adder_0/operator_B_stage_1_7/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_7/U2  ( .A(
        \adder_0/operator_B_stage_1_7/n3 ), .ZN(\adder_0/G1[7] ) );
  AND2_X1 \adder_0/operator_B_stage_1_7/U1  ( .A1(\adder_0/P0[13] ), .A2(
        \adder_0/P0[14] ), .ZN(\adder_0/P1[7] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_8/U3  ( .B1(\adder_0/G0[15] ), .B2(
        \adder_0/P0[16] ), .A(\adder_0/G0[16] ), .ZN(
        \adder_0/operator_B_stage_1_8/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_8/U2  ( .A(
        \adder_0/operator_B_stage_1_8/n3 ), .ZN(\adder_0/G1[8] ) );
  AND2_X1 \adder_0/operator_B_stage_1_8/U1  ( .A1(\adder_0/P0[15] ), .A2(
        \adder_0/P0[16] ), .ZN(\adder_0/P1[8] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_9/U3  ( .B1(\adder_0/G0[17] ), .B2(
        \adder_0/P0[18] ), .A(\adder_0/G0[18] ), .ZN(
        \adder_0/operator_B_stage_1_9/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_9/U2  ( .A(
        \adder_0/operator_B_stage_1_9/n3 ), .ZN(\adder_0/G1[9] ) );
  AND2_X1 \adder_0/operator_B_stage_1_9/U1  ( .A1(\adder_0/P0[17] ), .A2(
        \adder_0/P0[18] ), .ZN(\adder_0/P1[9] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_10/U3  ( .B1(\adder_0/G0[19] ), .B2(
        \adder_0/P0[20] ), .A(\adder_0/G0[20] ), .ZN(
        \adder_0/operator_B_stage_1_10/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_10/U2  ( .A(
        \adder_0/operator_B_stage_1_10/n3 ), .ZN(\adder_0/G1[10] ) );
  AND2_X1 \adder_0/operator_B_stage_1_10/U1  ( .A1(\adder_0/P0[19] ), .A2(
        \adder_0/P0[20] ), .ZN(\adder_0/P1[10] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_11/U3  ( .B1(\adder_0/G0[21] ), .B2(
        \adder_0/P0[22] ), .A(\adder_0/G0[22] ), .ZN(
        \adder_0/operator_B_stage_1_11/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_11/U2  ( .A(
        \adder_0/operator_B_stage_1_11/n3 ), .ZN(\adder_0/G1[11] ) );
  AND2_X1 \adder_0/operator_B_stage_1_11/U1  ( .A1(\adder_0/P0[21] ), .A2(
        \adder_0/P0[22] ), .ZN(\adder_0/P1[11] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_12/U3  ( .B1(\adder_0/G0[23] ), .B2(
        \adder_0/P0[24] ), .A(\adder_0/G0[24] ), .ZN(
        \adder_0/operator_B_stage_1_12/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_12/U2  ( .A(
        \adder_0/operator_B_stage_1_12/n3 ), .ZN(\adder_0/G1[12] ) );
  AND2_X1 \adder_0/operator_B_stage_1_12/U1  ( .A1(\adder_0/P0[23] ), .A2(
        \adder_0/P0[24] ), .ZN(\adder_0/P1[12] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_13/U3  ( .B1(\adder_0/G0[25] ), .B2(
        \adder_0/P0[26] ), .A(\adder_0/G0[26] ), .ZN(
        \adder_0/operator_B_stage_1_13/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_13/U2  ( .A(
        \adder_0/operator_B_stage_1_13/n3 ), .ZN(\adder_0/G1[13] ) );
  AND2_X1 \adder_0/operator_B_stage_1_13/U1  ( .A1(\adder_0/P0[25] ), .A2(
        \adder_0/P0[26] ), .ZN(\adder_0/P1[13] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_14/U3  ( .B1(\adder_0/G0[27] ), .B2(
        \adder_0/P0[28] ), .A(\adder_0/G0[28] ), .ZN(
        \adder_0/operator_B_stage_1_14/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_14/U2  ( .A(
        \adder_0/operator_B_stage_1_14/n3 ), .ZN(\adder_0/G1[14] ) );
  AND2_X1 \adder_0/operator_B_stage_1_14/U1  ( .A1(\adder_0/P0[27] ), .A2(
        \adder_0/P0[28] ), .ZN(\adder_0/P1[14] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_15/U3  ( .B1(\adder_0/G0[29] ), .B2(
        \adder_0/P0[30] ), .A(\adder_0/G0[30] ), .ZN(
        \adder_0/operator_B_stage_1_15/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_15/U2  ( .A(
        \adder_0/operator_B_stage_1_15/n3 ), .ZN(\adder_0/G1[15] ) );
  AND2_X1 \adder_0/operator_B_stage_1_15/U1  ( .A1(\adder_0/P0[29] ), .A2(
        \adder_0/P0[30] ), .ZN(\adder_0/P1[15] ) );
  AOI21_X1 \adder_0/operator_C_stage_2_1/U2  ( .B1(\adder_0/P1[1] ), .B2(
        \adder_0/G1[0] ), .A(\adder_0/G1[1] ), .ZN(
        \adder_0/operator_C_stage_2_1/n3 ) );
  INV_X1 \adder_0/operator_C_stage_2_1/U1  ( .A(
        \adder_0/operator_C_stage_2_1/n3 ), .ZN(\adder_0/G2[1] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_2/U3  ( .B1(\adder_0/G1[1] ), .B2(
        \adder_0/P1[2] ), .A(\adder_0/G1[2] ), .ZN(
        \adder_0/operator_B_stage_2_2/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_2/U2  ( .A(
        \adder_0/operator_B_stage_2_2/n3 ), .ZN(\adder_0/G2[2] ) );
  AND2_X1 \adder_0/operator_B_stage_2_2/U1  ( .A1(\adder_0/P1[1] ), .A2(
        \adder_0/P1[2] ), .ZN(\adder_0/P2[2] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_3/U3  ( .B1(\adder_0/G1[2] ), .B2(
        \adder_0/P1[3] ), .A(\adder_0/G1[3] ), .ZN(
        \adder_0/operator_B_stage_2_3/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_3/U2  ( .A(
        \adder_0/operator_B_stage_2_3/n3 ), .ZN(\adder_0/G2[3] ) );
  AND2_X1 \adder_0/operator_B_stage_2_3/U1  ( .A1(\adder_0/P1[2] ), .A2(
        \adder_0/P1[3] ), .ZN(\adder_0/P2[3] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_4/U3  ( .B1(\adder_0/G1[3] ), .B2(
        \adder_0/P1[4] ), .A(\adder_0/G1[4] ), .ZN(
        \adder_0/operator_B_stage_2_4/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_4/U2  ( .A(
        \adder_0/operator_B_stage_2_4/n3 ), .ZN(\adder_0/G2[4] ) );
  AND2_X1 \adder_0/operator_B_stage_2_4/U1  ( .A1(\adder_0/P1[3] ), .A2(
        \adder_0/P1[4] ), .ZN(\adder_0/P2[4] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_5/U3  ( .B1(\adder_0/G1[4] ), .B2(
        \adder_0/P1[5] ), .A(\adder_0/G1[5] ), .ZN(
        \adder_0/operator_B_stage_2_5/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_5/U2  ( .A(
        \adder_0/operator_B_stage_2_5/n3 ), .ZN(\adder_0/G2[5] ) );
  AND2_X1 \adder_0/operator_B_stage_2_5/U1  ( .A1(\adder_0/P1[4] ), .A2(
        \adder_0/P1[5] ), .ZN(\adder_0/P2[5] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_6/U3  ( .B1(\adder_0/G1[5] ), .B2(
        \adder_0/P1[6] ), .A(\adder_0/G1[6] ), .ZN(
        \adder_0/operator_B_stage_2_6/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_6/U2  ( .A(
        \adder_0/operator_B_stage_2_6/n3 ), .ZN(\adder_0/G2[6] ) );
  AND2_X1 \adder_0/operator_B_stage_2_6/U1  ( .A1(\adder_0/P1[5] ), .A2(
        \adder_0/P1[6] ), .ZN(\adder_0/P2[6] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_7/U3  ( .B1(\adder_0/G1[6] ), .B2(
        \adder_0/P1[7] ), .A(\adder_0/G1[7] ), .ZN(
        \adder_0/operator_B_stage_2_7/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_7/U2  ( .A(
        \adder_0/operator_B_stage_2_7/n3 ), .ZN(\adder_0/G2[7] ) );
  AND2_X1 \adder_0/operator_B_stage_2_7/U1  ( .A1(\adder_0/P1[6] ), .A2(
        \adder_0/P1[7] ), .ZN(\adder_0/P2[7] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_8/U3  ( .B1(\adder_0/G1[7] ), .B2(
        \adder_0/P1[8] ), .A(\adder_0/G1[8] ), .ZN(
        \adder_0/operator_B_stage_2_8/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_8/U2  ( .A(
        \adder_0/operator_B_stage_2_8/n3 ), .ZN(\adder_0/G2[8] ) );
  AND2_X1 \adder_0/operator_B_stage_2_8/U1  ( .A1(\adder_0/P1[7] ), .A2(
        \adder_0/P1[8] ), .ZN(\adder_0/P2[8] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_9/U3  ( .B1(\adder_0/G1[8] ), .B2(
        \adder_0/P1[9] ), .A(\adder_0/G1[9] ), .ZN(
        \adder_0/operator_B_stage_2_9/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_9/U2  ( .A(
        \adder_0/operator_B_stage_2_9/n3 ), .ZN(\adder_0/G2[9] ) );
  AND2_X1 \adder_0/operator_B_stage_2_9/U1  ( .A1(\adder_0/P1[8] ), .A2(
        \adder_0/P1[9] ), .ZN(\adder_0/P2[9] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_10/U3  ( .B1(\adder_0/G1[9] ), .B2(
        \adder_0/P1[10] ), .A(\adder_0/G1[10] ), .ZN(
        \adder_0/operator_B_stage_2_10/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_10/U2  ( .A(
        \adder_0/operator_B_stage_2_10/n3 ), .ZN(\adder_0/G2[10] ) );
  AND2_X1 \adder_0/operator_B_stage_2_10/U1  ( .A1(\adder_0/P1[9] ), .A2(
        \adder_0/P1[10] ), .ZN(\adder_0/P2[10] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_11/U3  ( .B1(\adder_0/G1[10] ), .B2(
        \adder_0/P1[11] ), .A(\adder_0/G1[11] ), .ZN(
        \adder_0/operator_B_stage_2_11/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_11/U2  ( .A(
        \adder_0/operator_B_stage_2_11/n3 ), .ZN(\adder_0/G2[11] ) );
  AND2_X1 \adder_0/operator_B_stage_2_11/U1  ( .A1(\adder_0/P1[10] ), .A2(
        \adder_0/P1[11] ), .ZN(\adder_0/P2[11] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_12/U3  ( .B1(\adder_0/G1[11] ), .B2(
        \adder_0/P1[12] ), .A(\adder_0/G1[12] ), .ZN(
        \adder_0/operator_B_stage_2_12/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_12/U2  ( .A(
        \adder_0/operator_B_stage_2_12/n3 ), .ZN(\adder_0/G2[12] ) );
  AND2_X1 \adder_0/operator_B_stage_2_12/U1  ( .A1(\adder_0/P1[11] ), .A2(
        \adder_0/P1[12] ), .ZN(\adder_0/P2[12] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_13/U3  ( .B1(\adder_0/G1[12] ), .B2(
        \adder_0/P1[13] ), .A(\adder_0/G1[13] ), .ZN(
        \adder_0/operator_B_stage_2_13/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_13/U2  ( .A(
        \adder_0/operator_B_stage_2_13/n3 ), .ZN(\adder_0/G2[13] ) );
  AND2_X1 \adder_0/operator_B_stage_2_13/U1  ( .A1(\adder_0/P1[12] ), .A2(
        \adder_0/P1[13] ), .ZN(\adder_0/P2[13] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_14/U3  ( .B1(\adder_0/G1[13] ), .B2(
        \adder_0/P1[14] ), .A(\adder_0/G1[14] ), .ZN(
        \adder_0/operator_B_stage_2_14/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_14/U2  ( .A(
        \adder_0/operator_B_stage_2_14/n3 ), .ZN(\adder_0/G2[14] ) );
  AND2_X1 \adder_0/operator_B_stage_2_14/U1  ( .A1(\adder_0/P1[13] ), .A2(
        \adder_0/P1[14] ), .ZN(\adder_0/P2[14] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_15/U3  ( .B1(\adder_0/G1[14] ), .B2(
        \adder_0/P1[15] ), .A(\adder_0/G1[15] ), .ZN(
        \adder_0/operator_B_stage_2_15/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_15/U2  ( .A(
        \adder_0/operator_B_stage_2_15/n3 ), .ZN(\adder_0/G2[15] ) );
  AND2_X1 \adder_0/operator_B_stage_2_15/U1  ( .A1(\adder_0/P1[14] ), .A2(
        \adder_0/P1[15] ), .ZN(\adder_0/P2[15] ) );
  AOI21_X1 \adder_0/operator_C_stage_3_2/U2  ( .B1(\adder_0/P2[2] ), .B2(
        \adder_0/G1[0] ), .A(\adder_0/G2[2] ), .ZN(
        \adder_0/operator_C_stage_3_2/n3 ) );
  INV_X1 \adder_0/operator_C_stage_3_2/U1  ( .A(
        \adder_0/operator_C_stage_3_2/n3 ), .ZN(\adder_0/G3[2] ) );
  AOI21_X1 \adder_0/operator_C_stage_3_3/U2  ( .B1(\adder_0/P2[3] ), .B2(
        \adder_0/G2[1] ), .A(\adder_0/G2[3] ), .ZN(
        \adder_0/operator_C_stage_3_3/n3 ) );
  INV_X1 \adder_0/operator_C_stage_3_3/U1  ( .A(
        \adder_0/operator_C_stage_3_3/n3 ), .ZN(\adder_0/G3[3] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_4/U3  ( .B1(\adder_0/G2[2] ), .B2(
        \adder_0/P2[4] ), .A(\adder_0/G2[4] ), .ZN(
        \adder_0/operator_B_stage_3_4/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_4/U2  ( .A(
        \adder_0/operator_B_stage_3_4/n3 ), .ZN(\adder_0/G3[4] ) );
  AND2_X1 \adder_0/operator_B_stage_3_4/U1  ( .A1(\adder_0/P2[2] ), .A2(
        \adder_0/P2[4] ), .ZN(\adder_0/P3[4] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_5/U3  ( .B1(\adder_0/G2[3] ), .B2(
        \adder_0/P2[5] ), .A(\adder_0/G2[5] ), .ZN(
        \adder_0/operator_B_stage_3_5/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_5/U2  ( .A(
        \adder_0/operator_B_stage_3_5/n3 ), .ZN(\adder_0/G3[5] ) );
  AND2_X1 \adder_0/operator_B_stage_3_5/U1  ( .A1(\adder_0/P2[3] ), .A2(
        \adder_0/P2[5] ), .ZN(\adder_0/P3[5] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_6/U3  ( .B1(\adder_0/G2[4] ), .B2(
        \adder_0/P2[6] ), .A(\adder_0/G2[6] ), .ZN(
        \adder_0/operator_B_stage_3_6/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_6/U2  ( .A(
        \adder_0/operator_B_stage_3_6/n3 ), .ZN(\adder_0/G3[6] ) );
  AND2_X1 \adder_0/operator_B_stage_3_6/U1  ( .A1(\adder_0/P2[4] ), .A2(
        \adder_0/P2[6] ), .ZN(\adder_0/P3[6] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_7/U3  ( .B1(\adder_0/G2[5] ), .B2(
        \adder_0/P2[7] ), .A(\adder_0/G2[7] ), .ZN(
        \adder_0/operator_B_stage_3_7/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_7/U2  ( .A(
        \adder_0/operator_B_stage_3_7/n3 ), .ZN(\adder_0/G3[7] ) );
  AND2_X1 \adder_0/operator_B_stage_3_7/U1  ( .A1(\adder_0/P2[5] ), .A2(
        \adder_0/P2[7] ), .ZN(\adder_0/P3[7] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_8/U3  ( .B1(\adder_0/G2[6] ), .B2(
        \adder_0/P2[8] ), .A(\adder_0/G2[8] ), .ZN(
        \adder_0/operator_B_stage_3_8/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_8/U2  ( .A(
        \adder_0/operator_B_stage_3_8/n3 ), .ZN(\adder_0/G3[8] ) );
  AND2_X1 \adder_0/operator_B_stage_3_8/U1  ( .A1(\adder_0/P2[6] ), .A2(
        \adder_0/P2[8] ), .ZN(\adder_0/P3[8] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_9/U3  ( .B1(\adder_0/G2[7] ), .B2(
        \adder_0/P2[9] ), .A(\adder_0/G2[9] ), .ZN(
        \adder_0/operator_B_stage_3_9/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_9/U2  ( .A(
        \adder_0/operator_B_stage_3_9/n3 ), .ZN(\adder_0/G3[9] ) );
  AND2_X1 \adder_0/operator_B_stage_3_9/U1  ( .A1(\adder_0/P2[7] ), .A2(
        \adder_0/P2[9] ), .ZN(\adder_0/P3[9] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_10/U3  ( .B1(\adder_0/G2[8] ), .B2(
        \adder_0/P2[10] ), .A(\adder_0/G2[10] ), .ZN(
        \adder_0/operator_B_stage_3_10/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_10/U2  ( .A(
        \adder_0/operator_B_stage_3_10/n3 ), .ZN(\adder_0/G3[10] ) );
  AND2_X1 \adder_0/operator_B_stage_3_10/U1  ( .A1(\adder_0/P2[8] ), .A2(
        \adder_0/P2[10] ), .ZN(\adder_0/P3[10] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_11/U3  ( .B1(\adder_0/G2[9] ), .B2(
        \adder_0/P2[11] ), .A(\adder_0/G2[11] ), .ZN(
        \adder_0/operator_B_stage_3_11/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_11/U2  ( .A(
        \adder_0/operator_B_stage_3_11/n3 ), .ZN(\adder_0/G3[11] ) );
  AND2_X1 \adder_0/operator_B_stage_3_11/U1  ( .A1(\adder_0/P2[9] ), .A2(
        \adder_0/P2[11] ), .ZN(\adder_0/P3[11] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_12/U3  ( .B1(\adder_0/G2[10] ), .B2(
        \adder_0/P2[12] ), .A(\adder_0/G2[12] ), .ZN(
        \adder_0/operator_B_stage_3_12/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_12/U2  ( .A(
        \adder_0/operator_B_stage_3_12/n3 ), .ZN(\adder_0/G3[12] ) );
  AND2_X1 \adder_0/operator_B_stage_3_12/U1  ( .A1(\adder_0/P2[10] ), .A2(
        \adder_0/P2[12] ), .ZN(\adder_0/P3[12] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_13/U3  ( .B1(\adder_0/G2[11] ), .B2(
        \adder_0/P2[13] ), .A(\adder_0/G2[13] ), .ZN(
        \adder_0/operator_B_stage_3_13/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_13/U2  ( .A(
        \adder_0/operator_B_stage_3_13/n3 ), .ZN(\adder_0/G3[13] ) );
  AND2_X1 \adder_0/operator_B_stage_3_13/U1  ( .A1(\adder_0/P2[11] ), .A2(
        \adder_0/P2[13] ), .ZN(\adder_0/P3[13] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_14/U3  ( .B1(\adder_0/G2[12] ), .B2(
        \adder_0/P2[14] ), .A(\adder_0/G2[14] ), .ZN(
        \adder_0/operator_B_stage_3_14/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_14/U2  ( .A(
        \adder_0/operator_B_stage_3_14/n3 ), .ZN(\adder_0/G3[14] ) );
  AND2_X1 \adder_0/operator_B_stage_3_14/U1  ( .A1(\adder_0/P2[12] ), .A2(
        \adder_0/P2[14] ), .ZN(\adder_0/P3[14] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_15/U3  ( .B1(\adder_0/G2[13] ), .B2(
        \adder_0/P2[15] ), .A(\adder_0/G2[15] ), .ZN(
        \adder_0/operator_B_stage_3_15/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_15/U2  ( .A(
        \adder_0/operator_B_stage_3_15/n3 ), .ZN(\adder_0/G3[15] ) );
  AND2_X1 \adder_0/operator_B_stage_3_15/U1  ( .A1(\adder_0/P2[13] ), .A2(
        \adder_0/P2[15] ), .ZN(\adder_0/P3[15] ) );
  AOI21_X1 \adder_0/operator_C_stage_4_4/U2  ( .B1(\adder_0/P3[4] ), .B2(
        \adder_0/G1[0] ), .A(\adder_0/G3[4] ), .ZN(
        \adder_0/operator_C_stage_4_4/n3 ) );
  INV_X1 \adder_0/operator_C_stage_4_4/U1  ( .A(
        \adder_0/operator_C_stage_4_4/n3 ), .ZN(\adder_0/G4[4] ) );
  AOI21_X1 \adder_0/operator_C_stage_4_5/U2  ( .B1(\adder_0/P3[5] ), .B2(
        \adder_0/G2[1] ), .A(\adder_0/G3[5] ), .ZN(
        \adder_0/operator_C_stage_4_5/n3 ) );
  INV_X1 \adder_0/operator_C_stage_4_5/U1  ( .A(
        \adder_0/operator_C_stage_4_5/n3 ), .ZN(\adder_0/G4[5] ) );
  AOI21_X1 \adder_0/operator_C_stage_4_6/U2  ( .B1(\adder_0/P3[6] ), .B2(
        \adder_0/G3[2] ), .A(\adder_0/G3[6] ), .ZN(
        \adder_0/operator_C_stage_4_6/n3 ) );
  INV_X1 \adder_0/operator_C_stage_4_6/U1  ( .A(
        \adder_0/operator_C_stage_4_6/n3 ), .ZN(\adder_0/G4[6] ) );
  AOI21_X1 \adder_0/operator_C_stage_4_7/U2  ( .B1(\adder_0/P3[7] ), .B2(
        \adder_0/G3[3] ), .A(\adder_0/G3[7] ), .ZN(
        \adder_0/operator_C_stage_4_7/n3 ) );
  INV_X1 \adder_0/operator_C_stage_4_7/U1  ( .A(
        \adder_0/operator_C_stage_4_7/n3 ), .ZN(\adder_0/G4[7] ) );
  AOI21_X1 \adder_0/operator_B_stage_4_8/U3  ( .B1(\adder_0/G3[4] ), .B2(
        \adder_0/P3[8] ), .A(\adder_0/G3[8] ), .ZN(
        \adder_0/operator_B_stage_4_8/n3 ) );
  INV_X1 \adder_0/operator_B_stage_4_8/U2  ( .A(
        \adder_0/operator_B_stage_4_8/n3 ), .ZN(\adder_0/G4[8] ) );
  AND2_X1 \adder_0/operator_B_stage_4_8/U1  ( .A1(\adder_0/P3[4] ), .A2(
        \adder_0/P3[8] ), .ZN(\adder_0/P4 [8]) );
  AOI21_X1 \adder_0/operator_B_stage_4_9/U3  ( .B1(\adder_0/G3[5] ), .B2(
        \adder_0/P3[9] ), .A(\adder_0/G3[9] ), .ZN(
        \adder_0/operator_B_stage_4_9/n3 ) );
  INV_X1 \adder_0/operator_B_stage_4_9/U2  ( .A(
        \adder_0/operator_B_stage_4_9/n3 ), .ZN(\adder_0/G4[9] ) );
  AND2_X1 \adder_0/operator_B_stage_4_9/U1  ( .A1(\adder_0/P3[5] ), .A2(
        \adder_0/P3[9] ), .ZN(\adder_0/P4 [9]) );
  AOI21_X1 \adder_0/operator_B_stage_4_10/U3  ( .B1(\adder_0/G3[6] ), .B2(
        \adder_0/P3[10] ), .A(\adder_0/G3[10] ), .ZN(
        \adder_0/operator_B_stage_4_10/n3 ) );
  INV_X1 \adder_0/operator_B_stage_4_10/U2  ( .A(
        \adder_0/operator_B_stage_4_10/n3 ), .ZN(\adder_0/G4[10] ) );
  AND2_X1 \adder_0/operator_B_stage_4_10/U1  ( .A1(\adder_0/P3[6] ), .A2(
        \adder_0/P3[10] ), .ZN(\adder_0/P4 [10]) );
  AOI21_X1 \adder_0/operator_B_stage_4_11/U3  ( .B1(\adder_0/G3[7] ), .B2(
        \adder_0/P3[11] ), .A(\adder_0/G3[11] ), .ZN(
        \adder_0/operator_B_stage_4_11/n3 ) );
  INV_X1 \adder_0/operator_B_stage_4_11/U2  ( .A(
        \adder_0/operator_B_stage_4_11/n3 ), .ZN(\adder_0/G4[11] ) );
  AND2_X1 \adder_0/operator_B_stage_4_11/U1  ( .A1(\adder_0/P3[7] ), .A2(
        \adder_0/P3[11] ), .ZN(\adder_0/P4 [11]) );
  AOI21_X1 \adder_0/operator_B_stage_4_12/U3  ( .B1(\adder_0/G3[8] ), .B2(
        \adder_0/P3[12] ), .A(\adder_0/G3[12] ), .ZN(
        \adder_0/operator_B_stage_4_12/n3 ) );
  INV_X1 \adder_0/operator_B_stage_4_12/U2  ( .A(
        \adder_0/operator_B_stage_4_12/n3 ), .ZN(\adder_0/G4[12] ) );
  AND2_X1 \adder_0/operator_B_stage_4_12/U1  ( .A1(\adder_0/P3[8] ), .A2(
        \adder_0/P3[12] ), .ZN(\adder_0/P4 [12]) );
  AOI21_X1 \adder_0/operator_B_stage_4_13/U3  ( .B1(\adder_0/G3[9] ), .B2(
        \adder_0/P3[13] ), .A(\adder_0/G3[13] ), .ZN(
        \adder_0/operator_B_stage_4_13/n3 ) );
  INV_X1 \adder_0/operator_B_stage_4_13/U2  ( .A(
        \adder_0/operator_B_stage_4_13/n3 ), .ZN(\adder_0/G4[13] ) );
  AND2_X1 \adder_0/operator_B_stage_4_13/U1  ( .A1(\adder_0/P3[9] ), .A2(
        \adder_0/P3[13] ), .ZN(\adder_0/P4 [13]) );
  AOI21_X1 \adder_0/operator_B_stage_4_14/U3  ( .B1(\adder_0/G3[10] ), .B2(
        \adder_0/P3[14] ), .A(\adder_0/G3[14] ), .ZN(
        \adder_0/operator_B_stage_4_14/n3 ) );
  INV_X1 \adder_0/operator_B_stage_4_14/U2  ( .A(
        \adder_0/operator_B_stage_4_14/n3 ), .ZN(\adder_0/G4[14] ) );
  AND2_X1 \adder_0/operator_B_stage_4_14/U1  ( .A1(\adder_0/P3[10] ), .A2(
        \adder_0/P3[14] ), .ZN(\adder_0/P4 [14]) );
  AOI21_X1 \adder_0/operator_B_stage_4_15/U3  ( .B1(\adder_0/G3[11] ), .B2(
        \adder_0/P3[15] ), .A(\adder_0/G3[15] ), .ZN(
        \adder_0/operator_B_stage_4_15/n3 ) );
  INV_X1 \adder_0/operator_B_stage_4_15/U2  ( .A(
        \adder_0/operator_B_stage_4_15/n3 ), .ZN(\adder_0/G4[15] ) );
  AND2_X1 \adder_0/operator_B_stage_4_15/U1  ( .A1(\adder_0/P3[11] ), .A2(
        \adder_0/P3[15] ), .ZN(\adder_0/P4 [15]) );
  AOI21_X1 \adder_0/operator_C_stage_5_8/U2  ( .B1(\adder_0/P4 [8]), .B2(
        \adder_0/G1[0] ), .A(\adder_0/G4[8] ), .ZN(
        \adder_0/operator_C_stage_5_8/n3 ) );
  INV_X1 \adder_0/operator_C_stage_5_8/U1  ( .A(
        \adder_0/operator_C_stage_5_8/n3 ), .ZN(\adder_0/G5[8] ) );
  AOI21_X1 \adder_0/operator_C_stage_5_9/U2  ( .B1(\adder_0/P4 [9]), .B2(
        \adder_0/G2[1] ), .A(\adder_0/G4[9] ), .ZN(
        \adder_0/operator_C_stage_5_9/n3 ) );
  INV_X1 \adder_0/operator_C_stage_5_9/U1  ( .A(
        \adder_0/operator_C_stage_5_9/n3 ), .ZN(\adder_0/G5[9] ) );
  AOI21_X1 \adder_0/operator_C_stage_5_10/U2  ( .B1(\adder_0/P4 [10]), .B2(
        \adder_0/G3[2] ), .A(\adder_0/G4[10] ), .ZN(
        \adder_0/operator_C_stage_5_10/n3 ) );
  INV_X1 \adder_0/operator_C_stage_5_10/U1  ( .A(
        \adder_0/operator_C_stage_5_10/n3 ), .ZN(\adder_0/G5[10] ) );
  AOI21_X1 \adder_0/operator_C_stage_5_11/U2  ( .B1(\adder_0/P4 [11]), .B2(
        \adder_0/G3[3] ), .A(\adder_0/G4[11] ), .ZN(
        \adder_0/operator_C_stage_5_11/n3 ) );
  INV_X1 \adder_0/operator_C_stage_5_11/U1  ( .A(
        \adder_0/operator_C_stage_5_11/n3 ), .ZN(\adder_0/G5[11] ) );
  AOI21_X1 \adder_0/operator_C_stage_5_12/U2  ( .B1(\adder_0/P4 [12]), .B2(
        \adder_0/G4[4] ), .A(\adder_0/G4[12] ), .ZN(
        \adder_0/operator_C_stage_5_12/n3 ) );
  INV_X1 \adder_0/operator_C_stage_5_12/U1  ( .A(
        \adder_0/operator_C_stage_5_12/n3 ), .ZN(\adder_0/G5[12] ) );
  AOI21_X1 \adder_0/operator_C_stage_5_13/U2  ( .B1(\adder_0/P4 [13]), .B2(
        \adder_0/G4[5] ), .A(\adder_0/G4[13] ), .ZN(
        \adder_0/operator_C_stage_5_13/n3 ) );
  INV_X1 \adder_0/operator_C_stage_5_13/U1  ( .A(
        \adder_0/operator_C_stage_5_13/n3 ), .ZN(\adder_0/G5[13] ) );
  AOI21_X1 \adder_0/operator_C_stage_5_14/U2  ( .B1(\adder_0/P4 [14]), .B2(
        \adder_0/G4[6] ), .A(\adder_0/G4[14] ), .ZN(
        \adder_0/operator_C_stage_5_14/n3 ) );
  INV_X1 \adder_0/operator_C_stage_5_14/U1  ( .A(
        \adder_0/operator_C_stage_5_14/n3 ), .ZN(\adder_0/G5[14] ) );
  AOI21_X1 \adder_0/operator_C_stage_5_15/U2  ( .B1(\adder_0/P4 [15]), .B2(
        \adder_0/G4[7] ), .A(\adder_0/G4[15] ), .ZN(
        \adder_0/operator_C_stage_5_15/n3 ) );
  INV_X1 \adder_0/operator_C_stage_5_15/U1  ( .A(
        \adder_0/operator_C_stage_5_15/n3 ), .ZN(\adder_0/G5[15] ) );
  AOI21_X1 \adder_0/operator_C_stage_6_0/U2  ( .B1(\adder_0/P0[1] ), .B2(
        \adder_0/G1[0] ), .A(\adder_0/G0[1] ), .ZN(
        \adder_0/operator_C_stage_6_0/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_0/U1  ( .A(
        \adder_0/operator_C_stage_6_0/n3 ), .ZN(\adder_0/G6_1 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_1/U2  ( .B1(\adder_0/P0[3] ), .B2(
        \adder_0/G2[1] ), .A(\adder_0/G0[3] ), .ZN(
        \adder_0/operator_C_stage_6_1/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_1/U1  ( .A(
        \adder_0/operator_C_stage_6_1/n3 ), .ZN(\adder_0/G6_3 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_2/U2  ( .B1(\adder_0/P0[5] ), .B2(
        \adder_0/G3[2] ), .A(\adder_0/G0[5] ), .ZN(
        \adder_0/operator_C_stage_6_2/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_2/U1  ( .A(
        \adder_0/operator_C_stage_6_2/n3 ), .ZN(\adder_0/G6_5 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_3/U2  ( .B1(\adder_0/P0[7] ), .B2(
        \adder_0/G3[3] ), .A(\adder_0/G0[7] ), .ZN(
        \adder_0/operator_C_stage_6_3/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_3/U1  ( .A(
        \adder_0/operator_C_stage_6_3/n3 ), .ZN(\adder_0/G6_7 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_4/U2  ( .B1(\adder_0/P0[9] ), .B2(
        \adder_0/G4[4] ), .A(\adder_0/G0[9] ), .ZN(
        \adder_0/operator_C_stage_6_4/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_4/U1  ( .A(
        \adder_0/operator_C_stage_6_4/n3 ), .ZN(\adder_0/G6_9 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_5/U2  ( .B1(\adder_0/P0[11] ), .B2(
        \adder_0/G4[5] ), .A(\adder_0/G0[11] ), .ZN(
        \adder_0/operator_C_stage_6_5/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_5/U1  ( .A(
        \adder_0/operator_C_stage_6_5/n3 ), .ZN(\adder_0/G6_11 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_6/U2  ( .B1(\adder_0/P0[13] ), .B2(
        \adder_0/G4[6] ), .A(\adder_0/G0[13] ), .ZN(
        \adder_0/operator_C_stage_6_6/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_6/U1  ( .A(
        \adder_0/operator_C_stage_6_6/n3 ), .ZN(\adder_0/G6_13 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_7/U2  ( .B1(\adder_0/P0[15] ), .B2(
        \adder_0/G4[7] ), .A(\adder_0/G0[15] ), .ZN(
        \adder_0/operator_C_stage_6_7/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_7/U1  ( .A(
        \adder_0/operator_C_stage_6_7/n3 ), .ZN(\adder_0/G6_15 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_8/U2  ( .B1(\adder_0/P0[17] ), .B2(
        \adder_0/G5[8] ), .A(\adder_0/G0[17] ), .ZN(
        \adder_0/operator_C_stage_6_8/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_8/U1  ( .A(
        \adder_0/operator_C_stage_6_8/n3 ), .ZN(\adder_0/G6_17 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_9/U2  ( .B1(\adder_0/P0[19] ), .B2(
        \adder_0/G5[9] ), .A(\adder_0/G0[19] ), .ZN(
        \adder_0/operator_C_stage_6_9/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_9/U1  ( .A(
        \adder_0/operator_C_stage_6_9/n3 ), .ZN(\adder_0/G6_19 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_10/U2  ( .B1(\adder_0/P0[21] ), .B2(
        \adder_0/G5[10] ), .A(\adder_0/G0[21] ), .ZN(
        \adder_0/operator_C_stage_6_10/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_10/U1  ( .A(
        \adder_0/operator_C_stage_6_10/n3 ), .ZN(\adder_0/G6_21 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_11/U2  ( .B1(\adder_0/P0[23] ), .B2(
        \adder_0/G5[11] ), .A(\adder_0/G0[23] ), .ZN(
        \adder_0/operator_C_stage_6_11/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_11/U1  ( .A(
        \adder_0/operator_C_stage_6_11/n3 ), .ZN(\adder_0/G6_23 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_12/U2  ( .B1(\adder_0/P0[25] ), .B2(
        \adder_0/G5[12] ), .A(\adder_0/G0[25] ), .ZN(
        \adder_0/operator_C_stage_6_12/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_12/U1  ( .A(
        \adder_0/operator_C_stage_6_12/n3 ), .ZN(\adder_0/G6_25 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_13/U2  ( .B1(\adder_0/P0[27] ), .B2(
        \adder_0/G5[13] ), .A(\adder_0/G0[27] ), .ZN(
        \adder_0/operator_C_stage_6_13/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_13/U1  ( .A(
        \adder_0/operator_C_stage_6_13/n3 ), .ZN(\adder_0/G6_27 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_14/U2  ( .B1(\adder_0/P0[29] ), .B2(
        \adder_0/G5[14] ), .A(\adder_0/G0[29] ), .ZN(
        \adder_0/operator_C_stage_6_14/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_14/U1  ( .A(
        \adder_0/operator_C_stage_6_14/n3 ), .ZN(\adder_0/G6_29_ ) );
  AOI21_X1 \adder_0/operator_C_stage_6_15/U2  ( .B1(\adder_0/P0[31] ), .B2(
        \adder_0/G5[15] ), .A(\adder_0/G0[31] ), .ZN(
        \adder_0/operator_C_stage_6_15/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_15/U1  ( .A(
        \adder_0/operator_C_stage_6_15/n3 ), .ZN(\adder_0/o_c ) );
  XOR2_X1 \adder_1/U32  ( .A(n1988), .B(\adder_1/P0[0] ), .Z(sum_ct[0]) );
  XOR2_X1 \adder_1/U31  ( .A(\adder_1/P0[10] ), .B(\adder_1/G6_9 ), .Z(
        SYNOPSYS_UNCONNECTED_23) );
  XOR2_X1 \adder_1/U30  ( .A(\adder_1/P0[11] ), .B(\adder_1/G4[5] ), .Z(
        SYNOPSYS_UNCONNECTED_22) );
  XOR2_X1 \adder_1/U29  ( .A(\adder_1/P0[12] ), .B(\adder_1/G6_11 ), .Z(
        SYNOPSYS_UNCONNECTED_21) );
  XOR2_X1 \adder_1/U28  ( .A(\adder_1/P0[13] ), .B(\adder_1/G4[6] ), .Z(
        SYNOPSYS_UNCONNECTED_20) );
  XOR2_X1 \adder_1/U27  ( .A(\adder_1/P0[14] ), .B(\adder_1/G6_13 ), .Z(
        SYNOPSYS_UNCONNECTED_19) );
  XOR2_X1 \adder_1/U26  ( .A(\adder_1/P0[15] ), .B(\adder_1/G4[7] ), .Z(
        SYNOPSYS_UNCONNECTED_18) );
  XOR2_X1 \adder_1/U25  ( .A(\adder_1/P0[16] ), .B(\adder_1/G6_15 ), .Z(
        SYNOPSYS_UNCONNECTED_17) );
  XOR2_X1 \adder_1/U24  ( .A(\adder_1/P0[17] ), .B(\adder_1/G5[8] ), .Z(
        SYNOPSYS_UNCONNECTED_16) );
  XOR2_X1 \adder_1/U23  ( .A(\adder_1/P0[18] ), .B(\adder_1/G6_17 ), .Z(
        SYNOPSYS_UNCONNECTED_15) );
  XOR2_X1 \adder_1/U22  ( .A(\adder_1/P0[19] ), .B(\adder_1/G5[9] ), .Z(
        SYNOPSYS_UNCONNECTED_14) );
  XOR2_X1 \adder_1/U21  ( .A(\adder_1/P0[1] ), .B(\adder_1/G1[0] ), .Z(
        sum_ct[1]) );
  XOR2_X1 \adder_1/U20  ( .A(\adder_1/P0[20] ), .B(\adder_1/G6_19 ), .Z(
        SYNOPSYS_UNCONNECTED_13) );
  XOR2_X1 \adder_1/U19  ( .A(\adder_1/P0[21] ), .B(\adder_1/G5[10] ), .Z(
        SYNOPSYS_UNCONNECTED_12) );
  XOR2_X1 \adder_1/U18  ( .A(\adder_1/P0[22] ), .B(\adder_1/G6_21 ), .Z(
        SYNOPSYS_UNCONNECTED_11) );
  XOR2_X1 \adder_1/U17  ( .A(\adder_1/P0[23] ), .B(\adder_1/G5[11] ), .Z(
        SYNOPSYS_UNCONNECTED_10) );
  XOR2_X1 \adder_1/U16  ( .A(\adder_1/P0[24] ), .B(\adder_1/G6_23 ), .Z(
        SYNOPSYS_UNCONNECTED_9) );
  XOR2_X1 \adder_1/U15  ( .A(\adder_1/P0[25] ), .B(\adder_1/G5[12] ), .Z(
        SYNOPSYS_UNCONNECTED_8) );
  XOR2_X1 \adder_1/U14  ( .A(\adder_1/P0[26] ), .B(\adder_1/G6_25 ), .Z(
        SYNOPSYS_UNCONNECTED_7) );
  XOR2_X1 \adder_1/U13  ( .A(\adder_1/P0[27] ), .B(\adder_1/G5[13] ), .Z(
        SYNOPSYS_UNCONNECTED_6) );
  XOR2_X1 \adder_1/U12  ( .A(\adder_1/P0[28] ), .B(\adder_1/G6_27 ), .Z(
        SYNOPSYS_UNCONNECTED_5) );
  XOR2_X1 \adder_1/U11  ( .A(\adder_1/P0[29] ), .B(\adder_1/G5[14] ), .Z(
        SYNOPSYS_UNCONNECTED_4) );
  XOR2_X1 \adder_1/U10  ( .A(\adder_1/P0[2] ), .B(\adder_1/G6_1 ), .Z(
        sum_ct[2]) );
  XOR2_X1 \adder_1/U9  ( .A(\adder_1/P0[30] ), .B(\adder_1/G6_29_ ), .Z(
        SYNOPSYS_UNCONNECTED_3) );
  XOR2_X1 \adder_1/U8  ( .A(\adder_1/P0[31] ), .B(\adder_1/G5[15] ), .Z(
        SYNOPSYS_UNCONNECTED_2) );
  XOR2_X1 \adder_1/U7  ( .A(\adder_1/P0[3] ), .B(\adder_1/G2[1] ), .Z(
        sum_ct[3]) );
  XOR2_X1 \adder_1/U6  ( .A(\adder_1/P0[4] ), .B(\adder_1/G6_3 ), .Z(sum_ct[4]) );
  XOR2_X1 \adder_1/U5  ( .A(\adder_1/P0[5] ), .B(\adder_1/G3[2] ), .Z(
        sum_ct[5]) );
  XOR2_X1 \adder_1/U4  ( .A(\adder_1/P0[6] ), .B(\adder_1/G6_5 ), .Z(
        SYNOPSYS_UNCONNECTED_27) );
  XOR2_X1 \adder_1/U3  ( .A(\adder_1/P0[7] ), .B(\adder_1/G3[3] ), .Z(
        SYNOPSYS_UNCONNECTED_26) );
  XOR2_X1 \adder_1/U2  ( .A(\adder_1/P0[8] ), .B(\adder_1/G6_7 ), .Z(
        SYNOPSYS_UNCONNECTED_25) );
  XOR2_X1 \adder_1/U1  ( .A(\adder_1/P0[9] ), .B(\adder_1/G4[4] ), .Z(
        SYNOPSYS_UNCONNECTED_24) );
  AND2_X1 \adder_1/operator_A_0/U2  ( .A1(n_1_net__0_), .A2(ct[0]), .ZN(
        \adder_1/G0[0] ) );
  XOR2_X1 \adder_1/operator_A_0/U1  ( .A(n_1_net__0_), .B(ct[0]), .Z(
        \adder_1/P0[0] ) );
  AND2_X1 \adder_1/operator_A_1/U2  ( .A1(n_1_net__1_), .A2(ct[1]), .ZN(
        \adder_1/G0[1] ) );
  XOR2_X1 \adder_1/operator_A_1/U1  ( .A(n_1_net__1_), .B(ct[1]), .Z(
        \adder_1/P0[1] ) );
  AND2_X1 \adder_1/operator_A_2/U2  ( .A1(n_1_net__2_), .A2(ct[2]), .ZN(
        \adder_1/G0[2] ) );
  XOR2_X1 \adder_1/operator_A_2/U1  ( .A(n_1_net__2_), .B(ct[2]), .Z(
        \adder_1/P0[2] ) );
  AND2_X1 \adder_1/operator_A_3/U2  ( .A1(n_1_net__3_), .A2(ct[3]), .ZN(
        \adder_1/G0[3] ) );
  XOR2_X1 \adder_1/operator_A_3/U1  ( .A(n_1_net__3_), .B(ct[3]), .Z(
        \adder_1/P0[3] ) );
  AND2_X1 \adder_1/operator_A_4/U2  ( .A1(n1988), .A2(ct[4]), .ZN(
        \adder_1/G0[4] ) );
  XOR2_X1 \adder_1/operator_A_4/U1  ( .A(n1988), .B(ct[4]), .Z(\adder_1/P0[4] ) );
  AND2_X1 \adder_1/operator_A_5/U2  ( .A1(n1988), .A2(ct[5]), .ZN(
        \adder_1/G0[5] ) );
  XOR2_X1 \adder_1/operator_A_5/U1  ( .A(n1988), .B(ct[5]), .Z(\adder_1/P0[5] ) );
  AND2_X1 \adder_1/operator_A_6/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[6] ) );
  XOR2_X1 \adder_1/operator_A_6/U1  ( .A(n1988), .B(1'b0), .Z(\adder_1/P0[6] )
         );
  AND2_X1 \adder_1/operator_A_7/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[7] ) );
  XOR2_X1 \adder_1/operator_A_7/U1  ( .A(n1988), .B(1'b0), .Z(\adder_1/P0[7] )
         );
  AND2_X1 \adder_1/operator_A_8/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[8] ) );
  XOR2_X1 \adder_1/operator_A_8/U1  ( .A(n1988), .B(1'b0), .Z(\adder_1/P0[8] )
         );
  AND2_X1 \adder_1/operator_A_9/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[9] ) );
  XOR2_X1 \adder_1/operator_A_9/U1  ( .A(n1988), .B(1'b0), .Z(\adder_1/P0[9] )
         );
  AND2_X1 \adder_1/operator_A_10/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[10] ) );
  XOR2_X1 \adder_1/operator_A_10/U1  ( .A(n1988), .B(1'b0), .Z(
        \adder_1/P0[10] ) );
  AND2_X1 \adder_1/operator_A_11/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[11] ) );
  XOR2_X1 \adder_1/operator_A_11/U1  ( .A(n1988), .B(1'b0), .Z(
        \adder_1/P0[11] ) );
  AND2_X1 \adder_1/operator_A_12/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[12] ) );
  XOR2_X1 \adder_1/operator_A_12/U1  ( .A(n1988), .B(1'b0), .Z(
        \adder_1/P0[12] ) );
  AND2_X1 \adder_1/operator_A_13/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[13] ) );
  XOR2_X1 \adder_1/operator_A_13/U1  ( .A(n1988), .B(1'b0), .Z(
        \adder_1/P0[13] ) );
  AND2_X1 \adder_1/operator_A_14/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[14] ) );
  XOR2_X1 \adder_1/operator_A_14/U1  ( .A(n1988), .B(1'b0), .Z(
        \adder_1/P0[14] ) );
  AND2_X1 \adder_1/operator_A_15/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[15] ) );
  XOR2_X1 \adder_1/operator_A_15/U1  ( .A(n1988), .B(1'b0), .Z(
        \adder_1/P0[15] ) );
  AND2_X1 \adder_1/operator_A_16/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[16] ) );
  XOR2_X1 \adder_1/operator_A_16/U1  ( .A(n1988), .B(1'b0), .Z(
        \adder_1/P0[16] ) );
  AND2_X1 \adder_1/operator_A_17/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[17] ) );
  XOR2_X1 \adder_1/operator_A_17/U1  ( .A(n1988), .B(1'b0), .Z(
        \adder_1/P0[17] ) );
  AND2_X1 \adder_1/operator_A_18/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[18] ) );
  XOR2_X1 \adder_1/operator_A_18/U1  ( .A(n1988), .B(1'b0), .Z(
        \adder_1/P0[18] ) );
  AND2_X1 \adder_1/operator_A_19/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[19] ) );
  XOR2_X1 \adder_1/operator_A_19/U1  ( .A(n1988), .B(1'b0), .Z(
        \adder_1/P0[19] ) );
  AND2_X1 \adder_1/operator_A_20/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[20] ) );
  XOR2_X1 \adder_1/operator_A_20/U1  ( .A(n1988), .B(1'b0), .Z(
        \adder_1/P0[20] ) );
  AND2_X1 \adder_1/operator_A_21/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[21] ) );
  XOR2_X1 \adder_1/operator_A_21/U1  ( .A(n1988), .B(1'b0), .Z(
        \adder_1/P0[21] ) );
  AND2_X1 \adder_1/operator_A_22/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[22] ) );
  XOR2_X1 \adder_1/operator_A_22/U1  ( .A(n1988), .B(1'b0), .Z(
        \adder_1/P0[22] ) );
  AND2_X1 \adder_1/operator_A_23/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[23] ) );
  XOR2_X1 \adder_1/operator_A_23/U1  ( .A(n1988), .B(1'b0), .Z(
        \adder_1/P0[23] ) );
  AND2_X1 \adder_1/operator_A_24/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[24] ) );
  XOR2_X1 \adder_1/operator_A_24/U1  ( .A(n1988), .B(1'b0), .Z(
        \adder_1/P0[24] ) );
  AND2_X1 \adder_1/operator_A_25/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[25] ) );
  XOR2_X1 \adder_1/operator_A_25/U1  ( .A(n1988), .B(1'b0), .Z(
        \adder_1/P0[25] ) );
  AND2_X1 \adder_1/operator_A_26/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[26] ) );
  XOR2_X1 \adder_1/operator_A_26/U1  ( .A(n1988), .B(1'b0), .Z(
        \adder_1/P0[26] ) );
  AND2_X1 \adder_1/operator_A_27/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[27] ) );
  XOR2_X1 \adder_1/operator_A_27/U1  ( .A(n1988), .B(1'b0), .Z(
        \adder_1/P0[27] ) );
  AND2_X1 \adder_1/operator_A_28/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[28] ) );
  XOR2_X1 \adder_1/operator_A_28/U1  ( .A(n1988), .B(1'b0), .Z(
        \adder_1/P0[28] ) );
  AND2_X1 \adder_1/operator_A_29/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[29] ) );
  XOR2_X1 \adder_1/operator_A_29/U1  ( .A(n1988), .B(1'b0), .Z(
        \adder_1/P0[29] ) );
  AND2_X1 \adder_1/operator_A_30/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[30] ) );
  XOR2_X1 \adder_1/operator_A_30/U1  ( .A(n1988), .B(1'b0), .Z(
        \adder_1/P0[30] ) );
  AND2_X1 \adder_1/operator_A_31/U2  ( .A1(n1988), .A2(1'b0), .ZN(
        \adder_1/G0[31] ) );
  XOR2_X1 \adder_1/operator_A_31/U1  ( .A(n1988), .B(1'b0), .Z(
        \adder_1/P0[31] ) );
  AOI21_X1 \adder_1/operator_C_stage_1_0/U2  ( .B1(\adder_1/P0[0] ), .B2(n1988), .A(\adder_1/G0[0] ), .ZN(\adder_1/operator_C_stage_1_0/n3 ) );
  INV_X1 \adder_1/operator_C_stage_1_0/U1  ( .A(
        \adder_1/operator_C_stage_1_0/n3 ), .ZN(\adder_1/G1[0] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_1/U3  ( .B1(\adder_1/G0[1] ), .B2(
        \adder_1/P0[2] ), .A(\adder_1/G0[2] ), .ZN(
        \adder_1/operator_B_stage_1_1/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_1/U2  ( .A(
        \adder_1/operator_B_stage_1_1/n3 ), .ZN(\adder_1/G1[1] ) );
  AND2_X1 \adder_1/operator_B_stage_1_1/U1  ( .A1(\adder_1/P0[1] ), .A2(
        \adder_1/P0[2] ), .ZN(\adder_1/P1[1] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_2/U3  ( .B1(\adder_1/G0[3] ), .B2(
        \adder_1/P0[4] ), .A(\adder_1/G0[4] ), .ZN(
        \adder_1/operator_B_stage_1_2/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_2/U2  ( .A(
        \adder_1/operator_B_stage_1_2/n3 ), .ZN(\adder_1/G1[2] ) );
  AND2_X1 \adder_1/operator_B_stage_1_2/U1  ( .A1(\adder_1/P0[3] ), .A2(
        \adder_1/P0[4] ), .ZN(\adder_1/P1[2] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_3/U3  ( .B1(\adder_1/G0[5] ), .B2(
        \adder_1/P0[6] ), .A(\adder_1/G0[6] ), .ZN(
        \adder_1/operator_B_stage_1_3/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_3/U2  ( .A(
        \adder_1/operator_B_stage_1_3/n3 ), .ZN(\adder_1/G1[3] ) );
  AND2_X1 \adder_1/operator_B_stage_1_3/U1  ( .A1(\adder_1/P0[5] ), .A2(
        \adder_1/P0[6] ), .ZN(\adder_1/P1[3] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_4/U3  ( .B1(\adder_1/G0[7] ), .B2(
        \adder_1/P0[8] ), .A(\adder_1/G0[8] ), .ZN(
        \adder_1/operator_B_stage_1_4/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_4/U2  ( .A(
        \adder_1/operator_B_stage_1_4/n3 ), .ZN(\adder_1/G1[4] ) );
  AND2_X1 \adder_1/operator_B_stage_1_4/U1  ( .A1(\adder_1/P0[7] ), .A2(
        \adder_1/P0[8] ), .ZN(\adder_1/P1[4] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_5/U3  ( .B1(\adder_1/G0[9] ), .B2(
        \adder_1/P0[10] ), .A(\adder_1/G0[10] ), .ZN(
        \adder_1/operator_B_stage_1_5/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_5/U2  ( .A(
        \adder_1/operator_B_stage_1_5/n3 ), .ZN(\adder_1/G1[5] ) );
  AND2_X1 \adder_1/operator_B_stage_1_5/U1  ( .A1(\adder_1/P0[9] ), .A2(
        \adder_1/P0[10] ), .ZN(\adder_1/P1[5] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_6/U3  ( .B1(\adder_1/G0[11] ), .B2(
        \adder_1/P0[12] ), .A(\adder_1/G0[12] ), .ZN(
        \adder_1/operator_B_stage_1_6/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_6/U2  ( .A(
        \adder_1/operator_B_stage_1_6/n3 ), .ZN(\adder_1/G1[6] ) );
  AND2_X1 \adder_1/operator_B_stage_1_6/U1  ( .A1(\adder_1/P0[11] ), .A2(
        \adder_1/P0[12] ), .ZN(\adder_1/P1[6] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_7/U3  ( .B1(\adder_1/G0[13] ), .B2(
        \adder_1/P0[14] ), .A(\adder_1/G0[14] ), .ZN(
        \adder_1/operator_B_stage_1_7/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_7/U2  ( .A(
        \adder_1/operator_B_stage_1_7/n3 ), .ZN(\adder_1/G1[7] ) );
  AND2_X1 \adder_1/operator_B_stage_1_7/U1  ( .A1(\adder_1/P0[13] ), .A2(
        \adder_1/P0[14] ), .ZN(\adder_1/P1[7] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_8/U3  ( .B1(\adder_1/G0[15] ), .B2(
        \adder_1/P0[16] ), .A(\adder_1/G0[16] ), .ZN(
        \adder_1/operator_B_stage_1_8/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_8/U2  ( .A(
        \adder_1/operator_B_stage_1_8/n3 ), .ZN(\adder_1/G1[8] ) );
  AND2_X1 \adder_1/operator_B_stage_1_8/U1  ( .A1(\adder_1/P0[15] ), .A2(
        \adder_1/P0[16] ), .ZN(\adder_1/P1[8] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_9/U3  ( .B1(\adder_1/G0[17] ), .B2(
        \adder_1/P0[18] ), .A(\adder_1/G0[18] ), .ZN(
        \adder_1/operator_B_stage_1_9/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_9/U2  ( .A(
        \adder_1/operator_B_stage_1_9/n3 ), .ZN(\adder_1/G1[9] ) );
  AND2_X1 \adder_1/operator_B_stage_1_9/U1  ( .A1(\adder_1/P0[17] ), .A2(
        \adder_1/P0[18] ), .ZN(\adder_1/P1[9] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_10/U3  ( .B1(\adder_1/G0[19] ), .B2(
        \adder_1/P0[20] ), .A(\adder_1/G0[20] ), .ZN(
        \adder_1/operator_B_stage_1_10/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_10/U2  ( .A(
        \adder_1/operator_B_stage_1_10/n3 ), .ZN(\adder_1/G1[10] ) );
  AND2_X1 \adder_1/operator_B_stage_1_10/U1  ( .A1(\adder_1/P0[19] ), .A2(
        \adder_1/P0[20] ), .ZN(\adder_1/P1[10] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_11/U3  ( .B1(\adder_1/G0[21] ), .B2(
        \adder_1/P0[22] ), .A(\adder_1/G0[22] ), .ZN(
        \adder_1/operator_B_stage_1_11/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_11/U2  ( .A(
        \adder_1/operator_B_stage_1_11/n3 ), .ZN(\adder_1/G1[11] ) );
  AND2_X1 \adder_1/operator_B_stage_1_11/U1  ( .A1(\adder_1/P0[21] ), .A2(
        \adder_1/P0[22] ), .ZN(\adder_1/P1[11] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_12/U3  ( .B1(\adder_1/G0[23] ), .B2(
        \adder_1/P0[24] ), .A(\adder_1/G0[24] ), .ZN(
        \adder_1/operator_B_stage_1_12/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_12/U2  ( .A(
        \adder_1/operator_B_stage_1_12/n3 ), .ZN(\adder_1/G1[12] ) );
  AND2_X1 \adder_1/operator_B_stage_1_12/U1  ( .A1(\adder_1/P0[23] ), .A2(
        \adder_1/P0[24] ), .ZN(\adder_1/P1[12] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_13/U3  ( .B1(\adder_1/G0[25] ), .B2(
        \adder_1/P0[26] ), .A(\adder_1/G0[26] ), .ZN(
        \adder_1/operator_B_stage_1_13/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_13/U2  ( .A(
        \adder_1/operator_B_stage_1_13/n3 ), .ZN(\adder_1/G1[13] ) );
  AND2_X1 \adder_1/operator_B_stage_1_13/U1  ( .A1(\adder_1/P0[25] ), .A2(
        \adder_1/P0[26] ), .ZN(\adder_1/P1[13] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_14/U3  ( .B1(\adder_1/G0[27] ), .B2(
        \adder_1/P0[28] ), .A(\adder_1/G0[28] ), .ZN(
        \adder_1/operator_B_stage_1_14/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_14/U2  ( .A(
        \adder_1/operator_B_stage_1_14/n3 ), .ZN(\adder_1/G1[14] ) );
  AND2_X1 \adder_1/operator_B_stage_1_14/U1  ( .A1(\adder_1/P0[27] ), .A2(
        \adder_1/P0[28] ), .ZN(\adder_1/P1[14] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_15/U3  ( .B1(\adder_1/G0[29] ), .B2(
        \adder_1/P0[30] ), .A(\adder_1/G0[30] ), .ZN(
        \adder_1/operator_B_stage_1_15/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_15/U2  ( .A(
        \adder_1/operator_B_stage_1_15/n3 ), .ZN(\adder_1/G1[15] ) );
  AND2_X1 \adder_1/operator_B_stage_1_15/U1  ( .A1(\adder_1/P0[29] ), .A2(
        \adder_1/P0[30] ), .ZN(\adder_1/P1[15] ) );
  AOI21_X1 \adder_1/operator_C_stage_2_1/U2  ( .B1(\adder_1/P1[1] ), .B2(
        \adder_1/G1[0] ), .A(\adder_1/G1[1] ), .ZN(
        \adder_1/operator_C_stage_2_1/n3 ) );
  INV_X1 \adder_1/operator_C_stage_2_1/U1  ( .A(
        \adder_1/operator_C_stage_2_1/n3 ), .ZN(\adder_1/G2[1] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_2/U3  ( .B1(\adder_1/G1[1] ), .B2(
        \adder_1/P1[2] ), .A(\adder_1/G1[2] ), .ZN(
        \adder_1/operator_B_stage_2_2/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_2/U2  ( .A(
        \adder_1/operator_B_stage_2_2/n3 ), .ZN(\adder_1/G2[2] ) );
  AND2_X1 \adder_1/operator_B_stage_2_2/U1  ( .A1(\adder_1/P1[1] ), .A2(
        \adder_1/P1[2] ), .ZN(\adder_1/P2[2] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_3/U3  ( .B1(\adder_1/G1[2] ), .B2(
        \adder_1/P1[3] ), .A(\adder_1/G1[3] ), .ZN(
        \adder_1/operator_B_stage_2_3/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_3/U2  ( .A(
        \adder_1/operator_B_stage_2_3/n3 ), .ZN(\adder_1/G2[3] ) );
  AND2_X1 \adder_1/operator_B_stage_2_3/U1  ( .A1(\adder_1/P1[2] ), .A2(
        \adder_1/P1[3] ), .ZN(\adder_1/P2[3] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_4/U3  ( .B1(\adder_1/G1[3] ), .B2(
        \adder_1/P1[4] ), .A(\adder_1/G1[4] ), .ZN(
        \adder_1/operator_B_stage_2_4/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_4/U2  ( .A(
        \adder_1/operator_B_stage_2_4/n3 ), .ZN(\adder_1/G2[4] ) );
  AND2_X1 \adder_1/operator_B_stage_2_4/U1  ( .A1(\adder_1/P1[3] ), .A2(
        \adder_1/P1[4] ), .ZN(\adder_1/P2[4] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_5/U3  ( .B1(\adder_1/G1[4] ), .B2(
        \adder_1/P1[5] ), .A(\adder_1/G1[5] ), .ZN(
        \adder_1/operator_B_stage_2_5/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_5/U2  ( .A(
        \adder_1/operator_B_stage_2_5/n3 ), .ZN(\adder_1/G2[5] ) );
  AND2_X1 \adder_1/operator_B_stage_2_5/U1  ( .A1(\adder_1/P1[4] ), .A2(
        \adder_1/P1[5] ), .ZN(\adder_1/P2[5] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_6/U3  ( .B1(\adder_1/G1[5] ), .B2(
        \adder_1/P1[6] ), .A(\adder_1/G1[6] ), .ZN(
        \adder_1/operator_B_stage_2_6/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_6/U2  ( .A(
        \adder_1/operator_B_stage_2_6/n3 ), .ZN(\adder_1/G2[6] ) );
  AND2_X1 \adder_1/operator_B_stage_2_6/U1  ( .A1(\adder_1/P1[5] ), .A2(
        \adder_1/P1[6] ), .ZN(\adder_1/P2[6] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_7/U3  ( .B1(\adder_1/G1[6] ), .B2(
        \adder_1/P1[7] ), .A(\adder_1/G1[7] ), .ZN(
        \adder_1/operator_B_stage_2_7/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_7/U2  ( .A(
        \adder_1/operator_B_stage_2_7/n3 ), .ZN(\adder_1/G2[7] ) );
  AND2_X1 \adder_1/operator_B_stage_2_7/U1  ( .A1(\adder_1/P1[6] ), .A2(
        \adder_1/P1[7] ), .ZN(\adder_1/P2[7] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_8/U3  ( .B1(\adder_1/G1[7] ), .B2(
        \adder_1/P1[8] ), .A(\adder_1/G1[8] ), .ZN(
        \adder_1/operator_B_stage_2_8/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_8/U2  ( .A(
        \adder_1/operator_B_stage_2_8/n3 ), .ZN(\adder_1/G2[8] ) );
  AND2_X1 \adder_1/operator_B_stage_2_8/U1  ( .A1(\adder_1/P1[7] ), .A2(
        \adder_1/P1[8] ), .ZN(\adder_1/P2[8] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_9/U3  ( .B1(\adder_1/G1[8] ), .B2(
        \adder_1/P1[9] ), .A(\adder_1/G1[9] ), .ZN(
        \adder_1/operator_B_stage_2_9/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_9/U2  ( .A(
        \adder_1/operator_B_stage_2_9/n3 ), .ZN(\adder_1/G2[9] ) );
  AND2_X1 \adder_1/operator_B_stage_2_9/U1  ( .A1(\adder_1/P1[8] ), .A2(
        \adder_1/P1[9] ), .ZN(\adder_1/P2[9] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_10/U3  ( .B1(\adder_1/G1[9] ), .B2(
        \adder_1/P1[10] ), .A(\adder_1/G1[10] ), .ZN(
        \adder_1/operator_B_stage_2_10/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_10/U2  ( .A(
        \adder_1/operator_B_stage_2_10/n3 ), .ZN(\adder_1/G2[10] ) );
  AND2_X1 \adder_1/operator_B_stage_2_10/U1  ( .A1(\adder_1/P1[9] ), .A2(
        \adder_1/P1[10] ), .ZN(\adder_1/P2[10] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_11/U3  ( .B1(\adder_1/G1[10] ), .B2(
        \adder_1/P1[11] ), .A(\adder_1/G1[11] ), .ZN(
        \adder_1/operator_B_stage_2_11/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_11/U2  ( .A(
        \adder_1/operator_B_stage_2_11/n3 ), .ZN(\adder_1/G2[11] ) );
  AND2_X1 \adder_1/operator_B_stage_2_11/U1  ( .A1(\adder_1/P1[10] ), .A2(
        \adder_1/P1[11] ), .ZN(\adder_1/P2[11] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_12/U3  ( .B1(\adder_1/G1[11] ), .B2(
        \adder_1/P1[12] ), .A(\adder_1/G1[12] ), .ZN(
        \adder_1/operator_B_stage_2_12/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_12/U2  ( .A(
        \adder_1/operator_B_stage_2_12/n3 ), .ZN(\adder_1/G2[12] ) );
  AND2_X1 \adder_1/operator_B_stage_2_12/U1  ( .A1(\adder_1/P1[11] ), .A2(
        \adder_1/P1[12] ), .ZN(\adder_1/P2[12] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_13/U3  ( .B1(\adder_1/G1[12] ), .B2(
        \adder_1/P1[13] ), .A(\adder_1/G1[13] ), .ZN(
        \adder_1/operator_B_stage_2_13/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_13/U2  ( .A(
        \adder_1/operator_B_stage_2_13/n3 ), .ZN(\adder_1/G2[13] ) );
  AND2_X1 \adder_1/operator_B_stage_2_13/U1  ( .A1(\adder_1/P1[12] ), .A2(
        \adder_1/P1[13] ), .ZN(\adder_1/P2[13] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_14/U3  ( .B1(\adder_1/G1[13] ), .B2(
        \adder_1/P1[14] ), .A(\adder_1/G1[14] ), .ZN(
        \adder_1/operator_B_stage_2_14/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_14/U2  ( .A(
        \adder_1/operator_B_stage_2_14/n3 ), .ZN(\adder_1/G2[14] ) );
  AND2_X1 \adder_1/operator_B_stage_2_14/U1  ( .A1(\adder_1/P1[13] ), .A2(
        \adder_1/P1[14] ), .ZN(\adder_1/P2[14] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_15/U3  ( .B1(\adder_1/G1[14] ), .B2(
        \adder_1/P1[15] ), .A(\adder_1/G1[15] ), .ZN(
        \adder_1/operator_B_stage_2_15/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_15/U2  ( .A(
        \adder_1/operator_B_stage_2_15/n3 ), .ZN(\adder_1/G2[15] ) );
  AND2_X1 \adder_1/operator_B_stage_2_15/U1  ( .A1(\adder_1/P1[14] ), .A2(
        \adder_1/P1[15] ), .ZN(\adder_1/P2[15] ) );
  AOI21_X1 \adder_1/operator_C_stage_3_2/U2  ( .B1(\adder_1/P2[2] ), .B2(
        \adder_1/G1[0] ), .A(\adder_1/G2[2] ), .ZN(
        \adder_1/operator_C_stage_3_2/n3 ) );
  INV_X1 \adder_1/operator_C_stage_3_2/U1  ( .A(
        \adder_1/operator_C_stage_3_2/n3 ), .ZN(\adder_1/G3[2] ) );
  AOI21_X1 \adder_1/operator_C_stage_3_3/U2  ( .B1(\adder_1/P2[3] ), .B2(
        \adder_1/G2[1] ), .A(\adder_1/G2[3] ), .ZN(
        \adder_1/operator_C_stage_3_3/n3 ) );
  INV_X1 \adder_1/operator_C_stage_3_3/U1  ( .A(
        \adder_1/operator_C_stage_3_3/n3 ), .ZN(\adder_1/G3[3] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_4/U3  ( .B1(\adder_1/G2[2] ), .B2(
        \adder_1/P2[4] ), .A(\adder_1/G2[4] ), .ZN(
        \adder_1/operator_B_stage_3_4/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_4/U2  ( .A(
        \adder_1/operator_B_stage_3_4/n3 ), .ZN(\adder_1/G3[4] ) );
  AND2_X1 \adder_1/operator_B_stage_3_4/U1  ( .A1(\adder_1/P2[2] ), .A2(
        \adder_1/P2[4] ), .ZN(\adder_1/P3[4] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_5/U3  ( .B1(\adder_1/G2[3] ), .B2(
        \adder_1/P2[5] ), .A(\adder_1/G2[5] ), .ZN(
        \adder_1/operator_B_stage_3_5/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_5/U2  ( .A(
        \adder_1/operator_B_stage_3_5/n3 ), .ZN(\adder_1/G3[5] ) );
  AND2_X1 \adder_1/operator_B_stage_3_5/U1  ( .A1(\adder_1/P2[3] ), .A2(
        \adder_1/P2[5] ), .ZN(\adder_1/P3[5] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_6/U3  ( .B1(\adder_1/G2[4] ), .B2(
        \adder_1/P2[6] ), .A(\adder_1/G2[6] ), .ZN(
        \adder_1/operator_B_stage_3_6/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_6/U2  ( .A(
        \adder_1/operator_B_stage_3_6/n3 ), .ZN(\adder_1/G3[6] ) );
  AND2_X1 \adder_1/operator_B_stage_3_6/U1  ( .A1(\adder_1/P2[4] ), .A2(
        \adder_1/P2[6] ), .ZN(\adder_1/P3[6] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_7/U3  ( .B1(\adder_1/G2[5] ), .B2(
        \adder_1/P2[7] ), .A(\adder_1/G2[7] ), .ZN(
        \adder_1/operator_B_stage_3_7/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_7/U2  ( .A(
        \adder_1/operator_B_stage_3_7/n3 ), .ZN(\adder_1/G3[7] ) );
  AND2_X1 \adder_1/operator_B_stage_3_7/U1  ( .A1(\adder_1/P2[5] ), .A2(
        \adder_1/P2[7] ), .ZN(\adder_1/P3[7] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_8/U3  ( .B1(\adder_1/G2[6] ), .B2(
        \adder_1/P2[8] ), .A(\adder_1/G2[8] ), .ZN(
        \adder_1/operator_B_stage_3_8/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_8/U2  ( .A(
        \adder_1/operator_B_stage_3_8/n3 ), .ZN(\adder_1/G3[8] ) );
  AND2_X1 \adder_1/operator_B_stage_3_8/U1  ( .A1(\adder_1/P2[6] ), .A2(
        \adder_1/P2[8] ), .ZN(\adder_1/P3[8] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_9/U3  ( .B1(\adder_1/G2[7] ), .B2(
        \adder_1/P2[9] ), .A(\adder_1/G2[9] ), .ZN(
        \adder_1/operator_B_stage_3_9/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_9/U2  ( .A(
        \adder_1/operator_B_stage_3_9/n3 ), .ZN(\adder_1/G3[9] ) );
  AND2_X1 \adder_1/operator_B_stage_3_9/U1  ( .A1(\adder_1/P2[7] ), .A2(
        \adder_1/P2[9] ), .ZN(\adder_1/P3[9] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_10/U3  ( .B1(\adder_1/G2[8] ), .B2(
        \adder_1/P2[10] ), .A(\adder_1/G2[10] ), .ZN(
        \adder_1/operator_B_stage_3_10/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_10/U2  ( .A(
        \adder_1/operator_B_stage_3_10/n3 ), .ZN(\adder_1/G3[10] ) );
  AND2_X1 \adder_1/operator_B_stage_3_10/U1  ( .A1(\adder_1/P2[8] ), .A2(
        \adder_1/P2[10] ), .ZN(\adder_1/P3[10] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_11/U3  ( .B1(\adder_1/G2[9] ), .B2(
        \adder_1/P2[11] ), .A(\adder_1/G2[11] ), .ZN(
        \adder_1/operator_B_stage_3_11/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_11/U2  ( .A(
        \adder_1/operator_B_stage_3_11/n3 ), .ZN(\adder_1/G3[11] ) );
  AND2_X1 \adder_1/operator_B_stage_3_11/U1  ( .A1(\adder_1/P2[9] ), .A2(
        \adder_1/P2[11] ), .ZN(\adder_1/P3[11] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_12/U3  ( .B1(\adder_1/G2[10] ), .B2(
        \adder_1/P2[12] ), .A(\adder_1/G2[12] ), .ZN(
        \adder_1/operator_B_stage_3_12/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_12/U2  ( .A(
        \adder_1/operator_B_stage_3_12/n3 ), .ZN(\adder_1/G3[12] ) );
  AND2_X1 \adder_1/operator_B_stage_3_12/U1  ( .A1(\adder_1/P2[10] ), .A2(
        \adder_1/P2[12] ), .ZN(\adder_1/P3[12] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_13/U3  ( .B1(\adder_1/G2[11] ), .B2(
        \adder_1/P2[13] ), .A(\adder_1/G2[13] ), .ZN(
        \adder_1/operator_B_stage_3_13/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_13/U2  ( .A(
        \adder_1/operator_B_stage_3_13/n3 ), .ZN(\adder_1/G3[13] ) );
  AND2_X1 \adder_1/operator_B_stage_3_13/U1  ( .A1(\adder_1/P2[11] ), .A2(
        \adder_1/P2[13] ), .ZN(\adder_1/P3[13] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_14/U3  ( .B1(\adder_1/G2[12] ), .B2(
        \adder_1/P2[14] ), .A(\adder_1/G2[14] ), .ZN(
        \adder_1/operator_B_stage_3_14/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_14/U2  ( .A(
        \adder_1/operator_B_stage_3_14/n3 ), .ZN(\adder_1/G3[14] ) );
  AND2_X1 \adder_1/operator_B_stage_3_14/U1  ( .A1(\adder_1/P2[12] ), .A2(
        \adder_1/P2[14] ), .ZN(\adder_1/P3[14] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_15/U3  ( .B1(\adder_1/G2[13] ), .B2(
        \adder_1/P2[15] ), .A(\adder_1/G2[15] ), .ZN(
        \adder_1/operator_B_stage_3_15/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_15/U2  ( .A(
        \adder_1/operator_B_stage_3_15/n3 ), .ZN(\adder_1/G3[15] ) );
  AND2_X1 \adder_1/operator_B_stage_3_15/U1  ( .A1(\adder_1/P2[13] ), .A2(
        \adder_1/P2[15] ), .ZN(\adder_1/P3[15] ) );
  AOI21_X1 \adder_1/operator_C_stage_4_4/U2  ( .B1(\adder_1/P3[4] ), .B2(
        \adder_1/G1[0] ), .A(\adder_1/G3[4] ), .ZN(
        \adder_1/operator_C_stage_4_4/n3 ) );
  INV_X1 \adder_1/operator_C_stage_4_4/U1  ( .A(
        \adder_1/operator_C_stage_4_4/n3 ), .ZN(\adder_1/G4[4] ) );
  AOI21_X1 \adder_1/operator_C_stage_4_5/U2  ( .B1(\adder_1/P3[5] ), .B2(
        \adder_1/G2[1] ), .A(\adder_1/G3[5] ), .ZN(
        \adder_1/operator_C_stage_4_5/n3 ) );
  INV_X1 \adder_1/operator_C_stage_4_5/U1  ( .A(
        \adder_1/operator_C_stage_4_5/n3 ), .ZN(\adder_1/G4[5] ) );
  AOI21_X1 \adder_1/operator_C_stage_4_6/U2  ( .B1(\adder_1/P3[6] ), .B2(
        \adder_1/G3[2] ), .A(\adder_1/G3[6] ), .ZN(
        \adder_1/operator_C_stage_4_6/n3 ) );
  INV_X1 \adder_1/operator_C_stage_4_6/U1  ( .A(
        \adder_1/operator_C_stage_4_6/n3 ), .ZN(\adder_1/G4[6] ) );
  AOI21_X1 \adder_1/operator_C_stage_4_7/U2  ( .B1(\adder_1/P3[7] ), .B2(
        \adder_1/G3[3] ), .A(\adder_1/G3[7] ), .ZN(
        \adder_1/operator_C_stage_4_7/n3 ) );
  INV_X1 \adder_1/operator_C_stage_4_7/U1  ( .A(
        \adder_1/operator_C_stage_4_7/n3 ), .ZN(\adder_1/G4[7] ) );
  AOI21_X1 \adder_1/operator_B_stage_4_8/U3  ( .B1(\adder_1/G3[4] ), .B2(
        \adder_1/P3[8] ), .A(\adder_1/G3[8] ), .ZN(
        \adder_1/operator_B_stage_4_8/n3 ) );
  INV_X1 \adder_1/operator_B_stage_4_8/U2  ( .A(
        \adder_1/operator_B_stage_4_8/n3 ), .ZN(\adder_1/G4[8] ) );
  AND2_X1 \adder_1/operator_B_stage_4_8/U1  ( .A1(\adder_1/P3[4] ), .A2(
        \adder_1/P3[8] ), .ZN(\adder_1/P4 [8]) );
  AOI21_X1 \adder_1/operator_B_stage_4_9/U3  ( .B1(\adder_1/G3[5] ), .B2(
        \adder_1/P3[9] ), .A(\adder_1/G3[9] ), .ZN(
        \adder_1/operator_B_stage_4_9/n3 ) );
  INV_X1 \adder_1/operator_B_stage_4_9/U2  ( .A(
        \adder_1/operator_B_stage_4_9/n3 ), .ZN(\adder_1/G4[9] ) );
  AND2_X1 \adder_1/operator_B_stage_4_9/U1  ( .A1(\adder_1/P3[5] ), .A2(
        \adder_1/P3[9] ), .ZN(\adder_1/P4 [9]) );
  AOI21_X1 \adder_1/operator_B_stage_4_10/U3  ( .B1(\adder_1/G3[6] ), .B2(
        \adder_1/P3[10] ), .A(\adder_1/G3[10] ), .ZN(
        \adder_1/operator_B_stage_4_10/n3 ) );
  INV_X1 \adder_1/operator_B_stage_4_10/U2  ( .A(
        \adder_1/operator_B_stage_4_10/n3 ), .ZN(\adder_1/G4[10] ) );
  AND2_X1 \adder_1/operator_B_stage_4_10/U1  ( .A1(\adder_1/P3[6] ), .A2(
        \adder_1/P3[10] ), .ZN(\adder_1/P4 [10]) );
  AOI21_X1 \adder_1/operator_B_stage_4_11/U3  ( .B1(\adder_1/G3[7] ), .B2(
        \adder_1/P3[11] ), .A(\adder_1/G3[11] ), .ZN(
        \adder_1/operator_B_stage_4_11/n3 ) );
  INV_X1 \adder_1/operator_B_stage_4_11/U2  ( .A(
        \adder_1/operator_B_stage_4_11/n3 ), .ZN(\adder_1/G4[11] ) );
  AND2_X1 \adder_1/operator_B_stage_4_11/U1  ( .A1(\adder_1/P3[7] ), .A2(
        \adder_1/P3[11] ), .ZN(\adder_1/P4 [11]) );
  AOI21_X1 \adder_1/operator_B_stage_4_12/U3  ( .B1(\adder_1/G3[8] ), .B2(
        \adder_1/P3[12] ), .A(\adder_1/G3[12] ), .ZN(
        \adder_1/operator_B_stage_4_12/n3 ) );
  INV_X1 \adder_1/operator_B_stage_4_12/U2  ( .A(
        \adder_1/operator_B_stage_4_12/n3 ), .ZN(\adder_1/G4[12] ) );
  AND2_X1 \adder_1/operator_B_stage_4_12/U1  ( .A1(\adder_1/P3[8] ), .A2(
        \adder_1/P3[12] ), .ZN(\adder_1/P4 [12]) );
  AOI21_X1 \adder_1/operator_B_stage_4_13/U3  ( .B1(\adder_1/G3[9] ), .B2(
        \adder_1/P3[13] ), .A(\adder_1/G3[13] ), .ZN(
        \adder_1/operator_B_stage_4_13/n3 ) );
  INV_X1 \adder_1/operator_B_stage_4_13/U2  ( .A(
        \adder_1/operator_B_stage_4_13/n3 ), .ZN(\adder_1/G4[13] ) );
  AND2_X1 \adder_1/operator_B_stage_4_13/U1  ( .A1(\adder_1/P3[9] ), .A2(
        \adder_1/P3[13] ), .ZN(\adder_1/P4 [13]) );
  AOI21_X1 \adder_1/operator_B_stage_4_14/U3  ( .B1(\adder_1/G3[10] ), .B2(
        \adder_1/P3[14] ), .A(\adder_1/G3[14] ), .ZN(
        \adder_1/operator_B_stage_4_14/n3 ) );
  INV_X1 \adder_1/operator_B_stage_4_14/U2  ( .A(
        \adder_1/operator_B_stage_4_14/n3 ), .ZN(\adder_1/G4[14] ) );
  AND2_X1 \adder_1/operator_B_stage_4_14/U1  ( .A1(\adder_1/P3[10] ), .A2(
        \adder_1/P3[14] ), .ZN(\adder_1/P4 [14]) );
  AOI21_X1 \adder_1/operator_B_stage_4_15/U3  ( .B1(\adder_1/G3[11] ), .B2(
        \adder_1/P3[15] ), .A(\adder_1/G3[15] ), .ZN(
        \adder_1/operator_B_stage_4_15/n3 ) );
  INV_X1 \adder_1/operator_B_stage_4_15/U2  ( .A(
        \adder_1/operator_B_stage_4_15/n3 ), .ZN(\adder_1/G4[15] ) );
  AND2_X1 \adder_1/operator_B_stage_4_15/U1  ( .A1(\adder_1/P3[11] ), .A2(
        \adder_1/P3[15] ), .ZN(\adder_1/P4 [15]) );
  AOI21_X1 \adder_1/operator_C_stage_5_8/U2  ( .B1(\adder_1/P4 [8]), .B2(
        \adder_1/G1[0] ), .A(\adder_1/G4[8] ), .ZN(
        \adder_1/operator_C_stage_5_8/n3 ) );
  INV_X1 \adder_1/operator_C_stage_5_8/U1  ( .A(
        \adder_1/operator_C_stage_5_8/n3 ), .ZN(\adder_1/G5[8] ) );
  AOI21_X1 \adder_1/operator_C_stage_5_9/U2  ( .B1(\adder_1/P4 [9]), .B2(
        \adder_1/G2[1] ), .A(\adder_1/G4[9] ), .ZN(
        \adder_1/operator_C_stage_5_9/n3 ) );
  INV_X1 \adder_1/operator_C_stage_5_9/U1  ( .A(
        \adder_1/operator_C_stage_5_9/n3 ), .ZN(\adder_1/G5[9] ) );
  AOI21_X1 \adder_1/operator_C_stage_5_10/U2  ( .B1(\adder_1/P4 [10]), .B2(
        \adder_1/G3[2] ), .A(\adder_1/G4[10] ), .ZN(
        \adder_1/operator_C_stage_5_10/n3 ) );
  INV_X1 \adder_1/operator_C_stage_5_10/U1  ( .A(
        \adder_1/operator_C_stage_5_10/n3 ), .ZN(\adder_1/G5[10] ) );
  AOI21_X1 \adder_1/operator_C_stage_5_11/U2  ( .B1(\adder_1/P4 [11]), .B2(
        \adder_1/G3[3] ), .A(\adder_1/G4[11] ), .ZN(
        \adder_1/operator_C_stage_5_11/n3 ) );
  INV_X1 \adder_1/operator_C_stage_5_11/U1  ( .A(
        \adder_1/operator_C_stage_5_11/n3 ), .ZN(\adder_1/G5[11] ) );
  AOI21_X1 \adder_1/operator_C_stage_5_12/U2  ( .B1(\adder_1/P4 [12]), .B2(
        \adder_1/G4[4] ), .A(\adder_1/G4[12] ), .ZN(
        \adder_1/operator_C_stage_5_12/n3 ) );
  INV_X1 \adder_1/operator_C_stage_5_12/U1  ( .A(
        \adder_1/operator_C_stage_5_12/n3 ), .ZN(\adder_1/G5[12] ) );
  AOI21_X1 \adder_1/operator_C_stage_5_13/U2  ( .B1(\adder_1/P4 [13]), .B2(
        \adder_1/G4[5] ), .A(\adder_1/G4[13] ), .ZN(
        \adder_1/operator_C_stage_5_13/n3 ) );
  INV_X1 \adder_1/operator_C_stage_5_13/U1  ( .A(
        \adder_1/operator_C_stage_5_13/n3 ), .ZN(\adder_1/G5[13] ) );
  AOI21_X1 \adder_1/operator_C_stage_5_14/U2  ( .B1(\adder_1/P4 [14]), .B2(
        \adder_1/G4[6] ), .A(\adder_1/G4[14] ), .ZN(
        \adder_1/operator_C_stage_5_14/n3 ) );
  INV_X1 \adder_1/operator_C_stage_5_14/U1  ( .A(
        \adder_1/operator_C_stage_5_14/n3 ), .ZN(\adder_1/G5[14] ) );
  AOI21_X1 \adder_1/operator_C_stage_5_15/U2  ( .B1(\adder_1/P4 [15]), .B2(
        \adder_1/G4[7] ), .A(\adder_1/G4[15] ), .ZN(
        \adder_1/operator_C_stage_5_15/n3 ) );
  INV_X1 \adder_1/operator_C_stage_5_15/U1  ( .A(
        \adder_1/operator_C_stage_5_15/n3 ), .ZN(\adder_1/G5[15] ) );
  AOI21_X1 \adder_1/operator_C_stage_6_0/U2  ( .B1(\adder_1/P0[1] ), .B2(
        \adder_1/G1[0] ), .A(\adder_1/G0[1] ), .ZN(
        \adder_1/operator_C_stage_6_0/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_0/U1  ( .A(
        \adder_1/operator_C_stage_6_0/n3 ), .ZN(\adder_1/G6_1 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_1/U2  ( .B1(\adder_1/P0[3] ), .B2(
        \adder_1/G2[1] ), .A(\adder_1/G0[3] ), .ZN(
        \adder_1/operator_C_stage_6_1/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_1/U1  ( .A(
        \adder_1/operator_C_stage_6_1/n3 ), .ZN(\adder_1/G6_3 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_2/U2  ( .B1(\adder_1/P0[5] ), .B2(
        \adder_1/G3[2] ), .A(\adder_1/G0[5] ), .ZN(
        \adder_1/operator_C_stage_6_2/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_2/U1  ( .A(
        \adder_1/operator_C_stage_6_2/n3 ), .ZN(\adder_1/G6_5 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_3/U2  ( .B1(\adder_1/P0[7] ), .B2(
        \adder_1/G3[3] ), .A(\adder_1/G0[7] ), .ZN(
        \adder_1/operator_C_stage_6_3/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_3/U1  ( .A(
        \adder_1/operator_C_stage_6_3/n3 ), .ZN(\adder_1/G6_7 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_4/U2  ( .B1(\adder_1/P0[9] ), .B2(
        \adder_1/G4[4] ), .A(\adder_1/G0[9] ), .ZN(
        \adder_1/operator_C_stage_6_4/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_4/U1  ( .A(
        \adder_1/operator_C_stage_6_4/n3 ), .ZN(\adder_1/G6_9 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_5/U2  ( .B1(\adder_1/P0[11] ), .B2(
        \adder_1/G4[5] ), .A(\adder_1/G0[11] ), .ZN(
        \adder_1/operator_C_stage_6_5/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_5/U1  ( .A(
        \adder_1/operator_C_stage_6_5/n3 ), .ZN(\adder_1/G6_11 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_6/U2  ( .B1(\adder_1/P0[13] ), .B2(
        \adder_1/G4[6] ), .A(\adder_1/G0[13] ), .ZN(
        \adder_1/operator_C_stage_6_6/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_6/U1  ( .A(
        \adder_1/operator_C_stage_6_6/n3 ), .ZN(\adder_1/G6_13 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_7/U2  ( .B1(\adder_1/P0[15] ), .B2(
        \adder_1/G4[7] ), .A(\adder_1/G0[15] ), .ZN(
        \adder_1/operator_C_stage_6_7/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_7/U1  ( .A(
        \adder_1/operator_C_stage_6_7/n3 ), .ZN(\adder_1/G6_15 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_8/U2  ( .B1(\adder_1/P0[17] ), .B2(
        \adder_1/G5[8] ), .A(\adder_1/G0[17] ), .ZN(
        \adder_1/operator_C_stage_6_8/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_8/U1  ( .A(
        \adder_1/operator_C_stage_6_8/n3 ), .ZN(\adder_1/G6_17 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_9/U2  ( .B1(\adder_1/P0[19] ), .B2(
        \adder_1/G5[9] ), .A(\adder_1/G0[19] ), .ZN(
        \adder_1/operator_C_stage_6_9/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_9/U1  ( .A(
        \adder_1/operator_C_stage_6_9/n3 ), .ZN(\adder_1/G6_19 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_10/U2  ( .B1(\adder_1/P0[21] ), .B2(
        \adder_1/G5[10] ), .A(\adder_1/G0[21] ), .ZN(
        \adder_1/operator_C_stage_6_10/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_10/U1  ( .A(
        \adder_1/operator_C_stage_6_10/n3 ), .ZN(\adder_1/G6_21 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_11/U2  ( .B1(\adder_1/P0[23] ), .B2(
        \adder_1/G5[11] ), .A(\adder_1/G0[23] ), .ZN(
        \adder_1/operator_C_stage_6_11/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_11/U1  ( .A(
        \adder_1/operator_C_stage_6_11/n3 ), .ZN(\adder_1/G6_23 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_12/U2  ( .B1(\adder_1/P0[25] ), .B2(
        \adder_1/G5[12] ), .A(\adder_1/G0[25] ), .ZN(
        \adder_1/operator_C_stage_6_12/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_12/U1  ( .A(
        \adder_1/operator_C_stage_6_12/n3 ), .ZN(\adder_1/G6_25 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_13/U2  ( .B1(\adder_1/P0[27] ), .B2(
        \adder_1/G5[13] ), .A(\adder_1/G0[27] ), .ZN(
        \adder_1/operator_C_stage_6_13/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_13/U1  ( .A(
        \adder_1/operator_C_stage_6_13/n3 ), .ZN(\adder_1/G6_27 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_14/U2  ( .B1(\adder_1/P0[29] ), .B2(
        \adder_1/G5[14] ), .A(\adder_1/G0[29] ), .ZN(
        \adder_1/operator_C_stage_6_14/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_14/U1  ( .A(
        \adder_1/operator_C_stage_6_14/n3 ), .ZN(\adder_1/G6_29_ ) );
  AOI21_X1 \adder_1/operator_C_stage_6_15/U2  ( .B1(\adder_1/P0[31] ), .B2(
        \adder_1/G5[15] ), .A(\adder_1/G0[31] ), .ZN(
        \adder_1/operator_C_stage_6_15/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_15/U1  ( .A(
        \adder_1/operator_C_stage_6_15/n3 ), .ZN(\adder_1/o_c ) );
  BUF_X1 \sra_198/U245  ( .A(PR_1[31]), .Z(N295) );
  INV_X1 \sra_198/U244  ( .A(PR_1[2]), .ZN(\sra_198/n257 ) );
  INV_X1 \sra_198/U243  ( .A(PR_1[27]), .ZN(\sra_198/n282 ) );
  INV_X1 \sra_198/U242  ( .A(PR_1[30]), .ZN(\sra_198/n285 ) );
  INV_X1 \sra_198/U241  ( .A(PR_1[3]), .ZN(\sra_198/n258 ) );
  INV_X1 \sra_198/U240  ( .A(PR_1[4]), .ZN(\sra_198/n259 ) );
  INV_X1 \sra_198/U239  ( .A(PR_1[5]), .ZN(\sra_198/n260 ) );
  INV_X1 \sra_198/U238  ( .A(PR_1[6]), .ZN(\sra_198/n261 ) );
  INV_X1 \sra_198/U237  ( .A(PR_1[18]), .ZN(\sra_198/n273 ) );
  INV_X1 \sra_198/U236  ( .A(PR_1[19]), .ZN(\sra_198/n274 ) );
  INV_X1 \sra_198/U235  ( .A(PR_1[14]), .ZN(\sra_198/n269 ) );
  INV_X1 \sra_198/U234  ( .A(PR_1[15]), .ZN(\sra_198/n270 ) );
  INV_X1 \sra_198/U233  ( .A(PR_1[11]), .ZN(\sra_198/n266 ) );
  INV_X1 \sra_198/U232  ( .A(PR_1[20]), .ZN(\sra_198/n275 ) );
  INV_X1 \sra_198/U231  ( .A(PR_1[16]), .ZN(\sra_198/n271 ) );
  INV_X1 \sra_198/U230  ( .A(PR_1[12]), .ZN(\sra_198/n267 ) );
  INV_X1 \sra_198/U229  ( .A(PR_1[21]), .ZN(\sra_198/n276 ) );
  INV_X1 \sra_198/U228  ( .A(PR_1[22]), .ZN(\sra_198/n277 ) );
  INV_X1 \sra_198/U227  ( .A(PR_1[23]), .ZN(\sra_198/n278 ) );
  INV_X1 \sra_198/U225  ( .A(PR_1[24]), .ZN(\sra_198/n279 ) );
  INV_X1 \sra_198/U224  ( .A(PR_1[25]), .ZN(\sra_198/n280 ) );
  INV_X1 \sra_198/U223  ( .A(PR_1[13]), .ZN(\sra_198/n268 ) );
  INV_X1 \sra_198/U222  ( .A(PR_1[17]), .ZN(\sra_198/n272 ) );
  INV_X1 \sra_198/U221  ( .A(PR_1[26]), .ZN(\sra_198/n281 ) );
  INV_X1 \sra_198/U220  ( .A(PR_1[28]), .ZN(\sra_198/n283 ) );
  INV_X1 \sra_198/U219  ( .A(PR_1[7]), .ZN(\sra_198/n262 ) );
  INV_X1 \sra_198/U218  ( .A(PR_1[8]), .ZN(\sra_198/n263 ) );
  INV_X1 \sra_198/U217  ( .A(PR_1[9]), .ZN(\sra_198/n264 ) );
  INV_X1 \sra_198/U216  ( .A(PR_1[10]), .ZN(\sra_198/n265 ) );
  INV_X1 \sra_198/U215  ( .A(PR_1[29]), .ZN(\sra_198/n284 ) );
  INV_X1 \sra_198/U214  ( .A(PR_1[31]), .ZN(\sra_198/n256 ) );
  INV_X1 \sra_198/U213  ( .A(ct_1[0]), .ZN(\sra_198/n255 ) );
  NAND2_X1 \sra_198/U212  ( .A1(ct_1[3]), .A2(PR_1[31]), .ZN(\sra_198/n163 )
         );
  INV_X1 \sra_198/U211  ( .A(ct_1[2]), .ZN(\sra_198/n241 ) );
  OAI221_X1 \sra_198/U210  ( .B1(\sra_198/n120 ), .B2(\sra_198/n257 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n258 ), .A(\sra_198/n212 ), .ZN(
        \sra_198/n200 ) );
  INV_X1 \sra_198/U209  ( .A(\sra_198/n201 ), .ZN(\sra_198/n222 ) );
  AOI21_X1 \sra_198/U208  ( .B1(\sra_198/n113 ), .B2(\sra_198/n200 ), .A(
        \sra_198/n222 ), .ZN(\sra_198/n199 ) );
  OAI221_X1 \sra_198/U207  ( .B1(\sra_198/n120 ), .B2(\sra_198/n258 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n259 ), .A(\sra_198/n161 ), .ZN(
        \sra_198/n155 ) );
  INV_X1 \sra_198/U205  ( .A(\sra_198/n156 ), .ZN(\sra_198/n221 ) );
  AOI21_X1 \sra_198/U204  ( .B1(\sra_198/n113 ), .B2(\sra_198/n155 ), .A(
        \sra_198/n221 ), .ZN(\sra_198/n154 ) );
  OAI221_X1 \sra_198/U203  ( .B1(\sra_198/n120 ), .B2(\sra_198/n259 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n260 ), .A(\sra_198/n134 ), .ZN(
        \sra_198/n129 ) );
  INV_X1 \sra_198/U202  ( .A(\sra_198/n130 ), .ZN(\sra_198/n220 ) );
  AOI21_X1 \sra_198/U201  ( .B1(\sra_198/n113 ), .B2(\sra_198/n129 ), .A(
        \sra_198/n220 ), .ZN(\sra_198/n128 ) );
  OAI221_X1 \sra_198/U200  ( .B1(\sra_198/n120 ), .B2(\sra_198/n260 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n261 ), .A(\sra_198/n125 ), .ZN(
        \sra_198/n114 ) );
  INV_X1 \sra_198/U199  ( .A(\sra_198/n115 ), .ZN(\sra_198/n219 ) );
  AOI21_X1 \sra_198/U198  ( .B1(\sra_198/n113 ), .B2(\sra_198/n114 ), .A(
        \sra_198/n219 ), .ZN(\sra_198/n111 ) );
  INV_X1 \sra_198/U197  ( .A(ct_1[3]), .ZN(\sra_198/n239 ) );
  NOR2_X1 \sra_198/U196  ( .A1(ct_1[4]), .A2(ct_1[5]), .ZN(\sra_198/n137 ) );
  NAND2_X1 \sra_198/U195  ( .A1(ct_1[5]), .A2(PR_1[31]), .ZN(\sra_198/n112 )
         );
  AOI22_X1 \sra_198/U194  ( .A1(PR_1[1]), .A2(\sra_198/n123 ), .B1(PR_1[0]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n212 ) );
  AOI22_X1 \sra_198/U193  ( .A1(PR_1[2]), .A2(\sra_198/n123 ), .B1(PR_1[1]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n161 ) );
  AOI22_X1 \sra_198/U192  ( .A1(PR_1[3]), .A2(\sra_198/n123 ), .B1(PR_1[2]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n134 ) );
  AOI22_X1 \sra_198/U191  ( .A1(PR_1[4]), .A2(\sra_198/n123 ), .B1(PR_1[3]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n125 ) );
  NAND2_X1 \sra_198/U190  ( .A1(ct_1[2]), .A2(\sra_198/n239 ), .ZN(
        \sra_198/n146 ) );
  NOR2_X1 \sra_198/U189  ( .A1(\sra_198/n147 ), .A2(ct_1[4]), .ZN(
        \sra_198/n113 ) );
  NAND2_X1 \sra_198/U188  ( .A1(\sra_198/n196 ), .A2(ct_1[2]), .ZN(
        \sra_198/n74 ) );
  AOI22_X1 \sra_198/U187  ( .A1(PR_1[5]), .A2(\sra_198/n123 ), .B1(PR_1[4]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n209 ) );
  OAI221_X1 \sra_198/U186  ( .B1(\sra_198/n120 ), .B2(\sra_198/n261 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n262 ), .A(\sra_198/n209 ), .ZN(
        \sra_198/n110 ) );
  AOI22_X1 \sra_198/U185  ( .A1(PR_1[6]), .A2(\sra_198/n123 ), .B1(PR_1[5]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n159 ) );
  OAI221_X1 \sra_198/U184  ( .B1(\sra_198/n120 ), .B2(\sra_198/n262 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n263 ), .A(\sra_198/n159 ), .ZN(
        \sra_198/n106 ) );
  AOI22_X1 \sra_198/U183  ( .A1(PR_1[7]), .A2(\sra_198/n123 ), .B1(PR_1[6]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n133 ) );
  OAI221_X1 \sra_198/U182  ( .B1(\sra_198/n120 ), .B2(\sra_198/n263 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n264 ), .A(\sra_198/n133 ), .ZN(
        \sra_198/n101 ) );
  AOI22_X1 \sra_198/U181  ( .A1(PR_1[8]), .A2(\sra_198/n123 ), .B1(PR_1[7]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n122 ) );
  OAI221_X1 \sra_198/U180  ( .B1(\sra_198/n120 ), .B2(\sra_198/n264 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n265 ), .A(\sra_198/n122 ), .ZN(
        \sra_198/n94 ) );
  AOI22_X1 \sra_198/U179  ( .A1(PR_1[21]), .A2(\sra_198/n123 ), .B1(PR_1[20]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n208 ) );
  OAI221_X1 \sra_198/U178  ( .B1(\sra_198/n120 ), .B2(\sra_198/n277 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n278 ), .A(\sra_198/n208 ), .ZN(
        \sra_198/n183 ) );
  AOI22_X1 \sra_198/U177  ( .A1(PR_1[23]), .A2(\sra_198/n123 ), .B1(PR_1[22]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n198 ) );
  OAI221_X1 \sra_198/U176  ( .B1(\sra_198/n120 ), .B2(\sra_198/n279 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n280 ), .A(\sra_198/n198 ), .ZN(
        \sra_198/n174 ) );
  AOI222_X1 \sra_198/U175  ( .A1(\sra_198/n124 ), .A2(PR_1[29]), .B1(
        \sra_198/n123 ), .B2(PR_1[30]), .C1(PR_1[31]), .C2(ct_1[1]), .ZN(
        \sra_198/n168 ) );
  OAI21_X1 \sra_198/U174  ( .B1(ct_1[5]), .B2(\sra_198/n199 ), .A(
        \sra_198/n112 ), .ZN(N264) );
  OAI21_X1 \sra_198/U173  ( .B1(ct_1[5]), .B2(\sra_198/n154 ), .A(
        \sra_198/n112 ), .ZN(N265) );
  OAI21_X1 \sra_198/U172  ( .B1(ct_1[5]), .B2(\sra_198/n128 ), .A(
        \sra_198/n112 ), .ZN(N266) );
  OAI21_X1 \sra_198/U171  ( .B1(ct_1[5]), .B2(\sra_198/n111 ), .A(
        \sra_198/n112 ), .ZN(N267) );
  OAI211_X1 \sra_198/U170  ( .C1(\sra_198/n244 ), .C2(\sra_198/n74 ), .A(
        \sra_198/n107 ), .B(\sra_198/n108 ), .ZN(N268) );
  OAI211_X1 \sra_198/U169  ( .C1(\sra_198/n245 ), .C2(\sra_198/n74 ), .A(
        \sra_198/n103 ), .B(\sra_198/n104 ), .ZN(N269) );
  OAI211_X1 \sra_198/U168  ( .C1(\sra_198/n252 ), .C2(\sra_198/n74 ), .A(
        \sra_198/n97 ), .B(\sra_198/n98 ), .ZN(N270) );
  OAI211_X1 \sra_198/U167  ( .C1(\sra_198/n249 ), .C2(\sra_198/n74 ), .A(
        \sra_198/n90 ), .B(\sra_198/n91 ), .ZN(N271) );
  OAI211_X1 \sra_198/U166  ( .C1(\sra_198/n243 ), .C2(\sra_198/n74 ), .A(
        \sra_198/n84 ), .B(\sra_198/n85 ), .ZN(N272) );
  OAI211_X1 \sra_198/U165  ( .C1(\sra_198/n246 ), .C2(\sra_198/n74 ), .A(
        \sra_198/n75 ), .B(\sra_198/n76 ), .ZN(N273) );
  OAI211_X1 \sra_198/U164  ( .C1(\sra_198/n253 ), .C2(\sra_198/n74 ), .A(
        \sra_198/n191 ), .B(\sra_198/n192 ), .ZN(N274) );
  OAI211_X1 \sra_198/U163  ( .C1(\sra_198/n250 ), .C2(\sra_198/n74 ), .A(
        \sra_198/n184 ), .B(\sra_198/n185 ), .ZN(N275) );
  OAI211_X1 \sra_198/U162  ( .C1(\sra_198/n254 ), .C2(\sra_198/n74 ), .A(
        \sra_198/n181 ), .B(\sra_198/n182 ), .ZN(N276) );
  OAI211_X1 \sra_198/U161  ( .C1(\sra_198/n247 ), .C2(\sra_198/n74 ), .A(
        \sra_198/n175 ), .B(\sra_198/n176 ), .ZN(N277) );
  OAI211_X1 \sra_198/U160  ( .C1(\sra_198/n251 ), .C2(\sra_198/n74 ), .A(
        \sra_198/n171 ), .B(\sra_198/n172 ), .ZN(N278) );
  OAI221_X1 \sra_198/U159  ( .B1(\sra_198/n250 ), .B2(\sra_198/n169 ), .C1(
        \sra_198/n248 ), .C2(\sra_198/n74 ), .A(\sra_198/n170 ), .ZN(N279) );
  OAI21_X1 \sra_198/U158  ( .B1(\sra_198/n235 ), .B2(\sra_198/n216 ), .A(
        \sra_198/n127 ), .ZN(N280) );
  OAI21_X1 \sra_198/U157  ( .B1(\sra_198/n158 ), .B2(\sra_198/n216 ), .A(
        \sra_198/n127 ), .ZN(N281) );
  OAI21_X1 \sra_198/U156  ( .B1(\sra_198/n132 ), .B2(\sra_198/n216 ), .A(
        \sra_198/n127 ), .ZN(N282) );
  OAI21_X1 \sra_198/U155  ( .B1(\sra_198/n117 ), .B2(\sra_198/n216 ), .A(
        \sra_198/n127 ), .ZN(N283) );
  OAI21_X1 \sra_198/U154  ( .B1(\sra_198/n234 ), .B2(\sra_198/n216 ), .A(
        \sra_198/n127 ), .ZN(N284) );
  OAI21_X1 \sra_198/U153  ( .B1(\sra_198/n233 ), .B2(\sra_198/n216 ), .A(
        \sra_198/n127 ), .ZN(N285) );
  OAI21_X1 \sra_198/U152  ( .B1(\sra_198/n232 ), .B2(\sra_198/n216 ), .A(
        \sra_198/n127 ), .ZN(N286) );
  OAI21_X1 \sra_198/U151  ( .B1(\sra_198/n93 ), .B2(\sra_198/n216 ), .A(
        \sra_198/n127 ), .ZN(N287) );
  OAI21_X1 \sra_198/U150  ( .B1(\sra_198/n87 ), .B2(\sra_198/n216 ), .A(
        \sra_198/n127 ), .ZN(N288) );
  OAI21_X1 \sra_198/U149  ( .B1(\sra_198/n80 ), .B2(\sra_198/n216 ), .A(
        \sra_198/n127 ), .ZN(N289) );
  OAI21_X1 \sra_198/U148  ( .B1(\sra_198/n140 ), .B2(\sra_198/n216 ), .A(
        \sra_198/n127 ), .ZN(N290) );
  OAI21_X1 \sra_198/U147  ( .B1(\sra_198/n139 ), .B2(\sra_198/n216 ), .A(
        \sra_198/n127 ), .ZN(N291) );
  OAI21_X1 \sra_198/U146  ( .B1(\sra_198/n138 ), .B2(\sra_198/n216 ), .A(
        \sra_198/n127 ), .ZN(N292) );
  INV_X1 \sra_198/U145  ( .A(\sra_198/n135 ), .ZN(N293) );
  OAI21_X1 \sra_198/U144  ( .B1(\sra_198/n126 ), .B2(\sra_198/n216 ), .A(
        \sra_198/n127 ), .ZN(N294) );
  AOI22_X1 \sra_198/U143  ( .A1(PR_1[27]), .A2(\sra_198/n123 ), .B1(PR_1[26]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n193 ) );
  OAI221_X1 \sra_198/U141  ( .B1(\sra_198/n120 ), .B2(\sra_198/n283 ), .C1(
        \sra_198/n284 ), .C2(\sra_198/n121 ), .A(\sra_198/n193 ), .ZN(
        \sra_198/n164 ) );
  AOI22_X1 \sra_198/U140  ( .A1(PR_1[24]), .A2(\sra_198/n123 ), .B1(PR_1[23]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n190 ) );
  OAI221_X1 \sra_198/U139  ( .B1(\sra_198/n120 ), .B2(\sra_198/n280 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n281 ), .A(\sra_198/n190 ), .ZN(
        \sra_198/n145 ) );
  AOI22_X1 \sra_198/U138  ( .A1(PR_1[9]), .A2(\sra_198/n123 ), .B1(PR_1[8]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n211 ) );
  OAI221_X1 \sra_198/U137  ( .B1(\sra_198/n120 ), .B2(\sra_198/n265 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n266 ), .A(\sra_198/n211 ), .ZN(
        \sra_198/n88 ) );
  AOI22_X1 \sra_198/U136  ( .A1(PR_1[10]), .A2(\sra_198/n123 ), .B1(PR_1[9]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n160 ) );
  OAI221_X1 \sra_198/U135  ( .B1(\sra_198/n120 ), .B2(\sra_198/n266 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n267 ), .A(\sra_198/n160 ), .ZN(
        \sra_198/n82 ) );
  AOI22_X1 \sra_198/U134  ( .A1(PR_1[11]), .A2(\sra_198/n123 ), .B1(PR_1[10]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n197 ) );
  OAI221_X1 \sra_198/U133  ( .B1(\sra_198/n120 ), .B2(\sra_198/n267 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n268 ), .A(\sra_198/n197 ), .ZN(
        \sra_198/n99 ) );
  AOI22_X1 \sra_198/U132  ( .A1(PR_1[12]), .A2(\sra_198/n123 ), .B1(PR_1[11]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n189 ) );
  OAI221_X1 \sra_198/U131  ( .B1(\sra_198/n120 ), .B2(\sra_198/n268 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n269 ), .A(\sra_198/n189 ), .ZN(
        \sra_198/n92 ) );
  AOI22_X1 \sra_198/U130  ( .A1(PR_1[17]), .A2(\sra_198/n123 ), .B1(PR_1[16]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n207 ) );
  OAI221_X1 \sra_198/U129  ( .B1(\sra_198/n120 ), .B2(\sra_198/n273 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n274 ), .A(\sra_198/n207 ), .ZN(
        \sra_198/n89 ) );
  AOI22_X1 \sra_198/U128  ( .A1(PR_1[19]), .A2(\sra_198/n123 ), .B1(PR_1[18]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n195 ) );
  OAI221_X1 \sra_198/U127  ( .B1(\sra_198/n120 ), .B2(\sra_198/n275 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n276 ), .A(\sra_198/n195 ), .ZN(
        \sra_198/n166 ) );
  AOI22_X1 \sra_198/U126  ( .A1(PR_1[25]), .A2(\sra_198/n123 ), .B1(PR_1[24]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n205 ) );
  OAI221_X1 \sra_198/U125  ( .B1(\sra_198/n120 ), .B2(\sra_198/n281 ), .C1(
        \sra_198/n282 ), .C2(\sra_198/n121 ), .A(\sra_198/n205 ), .ZN(
        \sra_198/n143 ) );
  AOI22_X1 \sra_198/U124  ( .A1(PR_1[26]), .A2(\sra_198/n123 ), .B1(PR_1[25]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n180 ) );
  OAI221_X1 \sra_198/U123  ( .B1(\sra_198/n120 ), .B2(\sra_198/n282 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n283 ), .A(\sra_198/n180 ), .ZN(
        \sra_198/n141 ) );
  AOI22_X1 \sra_198/U122  ( .A1(PR_1[22]), .A2(\sra_198/n123 ), .B1(PR_1[21]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n178 ) );
  OAI221_X1 \sra_198/U121  ( .B1(\sra_198/n120 ), .B2(\sra_198/n278 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n279 ), .A(\sra_198/n178 ), .ZN(
        \sra_198/n152 ) );
  AOI22_X1 \sra_198/U120  ( .A1(PR_1[28]), .A2(\sra_198/n123 ), .B1(PR_1[27]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n186 ) );
  OAI221_X1 \sra_198/U119  ( .B1(\sra_198/n284 ), .B2(\sra_198/n120 ), .C1(
        \sra_198/n285 ), .C2(\sra_198/n121 ), .A(\sra_198/n186 ), .ZN(
        \sra_198/n144 ) );
  NAND2_X1 \sra_198/U118  ( .A1(PR_1[31]), .A2(\sra_198/n216 ), .ZN(
        \sra_198/n127 ) );
  AOI22_X1 \sra_198/U117  ( .A1(PR_1[29]), .A2(\sra_198/n123 ), .B1(PR_1[28]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n206 ) );
  OAI221_X1 \sra_198/U116  ( .B1(\sra_198/n285 ), .B2(\sra_198/n120 ), .C1(
        \sra_198/n256 ), .C2(\sra_198/n121 ), .A(\sra_198/n206 ), .ZN(
        \sra_198/n142 ) );
  AOI22_X1 \sra_198/U114  ( .A1(PR_1[16]), .A2(\sra_198/n123 ), .B1(PR_1[15]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n187 ) );
  OAI221_X1 \sra_198/U113  ( .B1(\sra_198/n120 ), .B2(\sra_198/n272 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n273 ), .A(\sra_198/n187 ), .ZN(
        \sra_198/n95 ) );
  AOI22_X1 \sra_198/U112  ( .A1(PR_1[18]), .A2(\sra_198/n123 ), .B1(PR_1[17]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n177 ) );
  OAI221_X1 \sra_198/U111  ( .B1(\sra_198/n120 ), .B2(\sra_198/n274 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n275 ), .A(\sra_198/n177 ), .ZN(
        \sra_198/n83 ) );
  AOI22_X1 \sra_198/U110  ( .A1(PR_1[13]), .A2(\sra_198/n123 ), .B1(PR_1[12]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n210 ) );
  OAI221_X1 \sra_198/U109  ( .B1(\sra_198/n120 ), .B2(\sra_198/n269 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n270 ), .A(\sra_198/n210 ), .ZN(
        \sra_198/n86 ) );
  AOI22_X1 \sra_198/U108  ( .A1(PR_1[14]), .A2(\sra_198/n123 ), .B1(PR_1[13]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n179 ) );
  OAI221_X1 \sra_198/U107  ( .B1(\sra_198/n120 ), .B2(\sra_198/n270 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n271 ), .A(\sra_198/n179 ), .ZN(
        \sra_198/n78 ) );
  AOI22_X1 \sra_198/U105  ( .A1(PR_1[15]), .A2(\sra_198/n123 ), .B1(PR_1[14]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n194 ) );
  OAI221_X1 \sra_198/U104  ( .B1(\sra_198/n120 ), .B2(\sra_198/n271 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n272 ), .A(\sra_198/n194 ), .ZN(
        \sra_198/n102 ) );
  AOI22_X1 \sra_198/U103  ( .A1(PR_1[20]), .A2(\sra_198/n123 ), .B1(PR_1[19]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n188 ) );
  OAI221_X1 \sra_198/U102  ( .B1(\sra_198/n120 ), .B2(\sra_198/n276 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n277 ), .A(\sra_198/n188 ), .ZN(
        \sra_198/n96 ) );
  INV_X1 \sra_198/U101  ( .A(ct_1[4]), .ZN(\sra_198/n218 ) );
  AOI22_X1 \sra_198/U100  ( .A1(\sra_198/n119 ), .A2(\sra_198/n142 ), .B1(
        \sra_198/n118 ), .B2(\sra_198/n143 ), .ZN(\sra_198/n204 ) );
  OAI221_X1 \sra_198/U99  ( .B1(\sra_198/n243 ), .B2(\sra_198/n146 ), .C1(
        \sra_198/n244 ), .C2(\sra_198/n147 ), .A(\sra_198/n204 ), .ZN(
        \sra_198/n203 ) );
  INV_X1 \sra_198/U98  ( .A(\sra_198/n203 ), .ZN(\sra_198/n235 ) );
  NAND2_X1 \sra_198/U97  ( .A1(\sra_198/n196 ), .A2(\sra_198/n241 ), .ZN(
        \sra_198/n169 ) );
  INV_X1 \sra_198/U96  ( .A(\sra_198/n144 ), .ZN(\sra_198/n248 ) );
  INV_X1 \sra_198/U95  ( .A(\sra_198/n83 ), .ZN(\sra_198/n245 ) );
  INV_X1 \sra_198/U94  ( .A(\sra_198/n96 ), .ZN(\sra_198/n249 ) );
  INV_X1 \sra_198/U93  ( .A(\sra_198/n89 ), .ZN(\sra_198/n244 ) );
  INV_X1 \sra_198/U92  ( .A(\sra_198/n152 ), .ZN(\sra_198/n246 ) );
  INV_X1 \sra_198/U91  ( .A(\sra_198/n166 ), .ZN(\sra_198/n252 ) );
  INV_X1 \sra_198/U90  ( .A(\sra_198/n145 ), .ZN(\sra_198/n250 ) );
  INV_X1 \sra_198/U89  ( .A(\sra_198/n141 ), .ZN(\sra_198/n247 ) );
  INV_X1 \sra_198/U88  ( .A(\sra_198/n164 ), .ZN(\sra_198/n251 ) );
  INV_X1 \sra_198/U87  ( .A(\sra_198/n143 ), .ZN(\sra_198/n254 ) );
  INV_X1 \sra_198/U86  ( .A(\sra_198/n174 ), .ZN(\sra_198/n253 ) );
  INV_X1 \sra_198/U85  ( .A(\sra_198/n183 ), .ZN(\sra_198/n243 ) );
  INV_X1 \sra_198/U84  ( .A(\sra_198/n163 ), .ZN(\sra_198/n240 ) );
  INV_X1 \sra_198/U83  ( .A(\sra_198/n127 ), .ZN(\sra_198/n215 ) );
  AOI21_X1 \sra_198/U82  ( .B1(\sra_198/n136 ), .B2(\sra_198/n137 ), .A(
        \sra_198/n215 ), .ZN(\sra_198/n135 ) );
  INV_X1 \sra_198/U81  ( .A(\sra_198/n168 ), .ZN(\sra_198/n242 ) );
  NOR2_X1 \sra_198/U80  ( .A1(\sra_198/n216 ), .A2(\sra_198/n239 ), .ZN(
        \sra_198/n196 ) );
  AOI21_X1 \sra_198/U79  ( .B1(\sra_198/n149 ), .B2(\sra_198/n231 ), .A(
        \sra_198/n173 ), .ZN(\sra_198/n126 ) );
  AOI22_X1 \sra_198/U78  ( .A1(\sra_198/n81 ), .A2(\sra_198/n110 ), .B1(
        \sra_198/n214 ), .B2(\sra_198/n86 ), .ZN(\sra_198/n107 ) );
  AOI22_X1 \sra_198/U77  ( .A1(\sra_198/n81 ), .A2(\sra_198/n106 ), .B1(
        \sra_198/n214 ), .B2(\sra_198/n78 ), .ZN(\sra_198/n103 ) );
  AOI22_X1 \sra_198/U76  ( .A1(\sra_198/n81 ), .A2(\sra_198/n101 ), .B1(
        \sra_198/n214 ), .B2(\sra_198/n102 ), .ZN(\sra_198/n97 ) );
  AOI22_X1 \sra_198/U75  ( .A1(\sra_198/n81 ), .A2(\sra_198/n94 ), .B1(
        \sra_198/n214 ), .B2(\sra_198/n95 ), .ZN(\sra_198/n90 ) );
  AOI22_X1 \sra_198/U74  ( .A1(\sra_198/n81 ), .A2(\sra_198/n88 ), .B1(
        \sra_198/n214 ), .B2(\sra_198/n89 ), .ZN(\sra_198/n84 ) );
  AOI22_X1 \sra_198/U73  ( .A1(\sra_198/n81 ), .A2(\sra_198/n82 ), .B1(
        \sra_198/n214 ), .B2(\sra_198/n83 ), .ZN(\sra_198/n75 ) );
  AOI22_X1 \sra_198/U72  ( .A1(\sra_198/n81 ), .A2(\sra_198/n99 ), .B1(
        \sra_198/n214 ), .B2(\sra_198/n166 ), .ZN(\sra_198/n191 ) );
  AOI22_X1 \sra_198/U71  ( .A1(\sra_198/n81 ), .A2(\sra_198/n92 ), .B1(
        \sra_198/n214 ), .B2(\sra_198/n96 ), .ZN(\sra_198/n184 ) );
  AOI22_X1 \sra_198/U70  ( .A1(\sra_198/n81 ), .A2(\sra_198/n86 ), .B1(
        \sra_198/n214 ), .B2(\sra_198/n183 ), .ZN(\sra_198/n181 ) );
  AOI22_X1 \sra_198/U69  ( .A1(\sra_198/n81 ), .A2(\sra_198/n78 ), .B1(
        \sra_198/n214 ), .B2(\sra_198/n152 ), .ZN(\sra_198/n175 ) );
  AOI22_X1 \sra_198/U68  ( .A1(\sra_198/n81 ), .A2(\sra_198/n102 ), .B1(
        \sra_198/n214 ), .B2(\sra_198/n174 ), .ZN(\sra_198/n171 ) );
  AOI21_X1 \sra_198/U67  ( .B1(\sra_198/n144 ), .B2(\sra_198/n231 ), .A(
        \sra_198/n173 ), .ZN(\sra_198/n139 ) );
  AOI21_X1 \sra_198/U66  ( .B1(\sra_198/n142 ), .B2(\sra_198/n231 ), .A(
        \sra_198/n173 ), .ZN(\sra_198/n138 ) );
  INV_X1 \sra_198/U65  ( .A(\sra_198/n173 ), .ZN(\sra_198/n224 ) );
  OAI21_X1 \sra_198/U64  ( .B1(\sra_198/n168 ), .B2(\sra_198/n147 ), .A(
        \sra_198/n224 ), .ZN(\sra_198/n136 ) );
  AOI222_X1 \sra_198/U63  ( .A1(\sra_198/n88 ), .A2(\sra_198/n118 ), .B1(
        \sra_198/n86 ), .B2(\sra_198/n119 ), .C1(\sra_198/n110 ), .C2(
        \sra_198/n238 ), .ZN(\sra_198/n202 ) );
  AOI222_X1 \sra_198/U62  ( .A1(\sra_198/n82 ), .A2(\sra_198/n118 ), .B1(
        \sra_198/n78 ), .B2(\sra_198/n119 ), .C1(\sra_198/n106 ), .C2(
        \sra_198/n238 ), .ZN(\sra_198/n157 ) );
  AOI222_X1 \sra_198/U61  ( .A1(\sra_198/n99 ), .A2(\sra_198/n118 ), .B1(
        \sra_198/n102 ), .B2(\sra_198/n119 ), .C1(\sra_198/n101 ), .C2(
        \sra_198/n238 ), .ZN(\sra_198/n131 ) );
  AOI222_X1 \sra_198/U60  ( .A1(\sra_198/n92 ), .A2(\sra_198/n118 ), .B1(
        \sra_198/n95 ), .B2(\sra_198/n119 ), .C1(\sra_198/n94 ), .C2(
        \sra_198/n238 ), .ZN(\sra_198/n116 ) );
  NOR2_X1 \sra_198/U59  ( .A1(\sra_198/n163 ), .A2(\sra_198/n241 ), .ZN(
        \sra_198/n150 ) );
  NOR2_X1 \sra_198/U58  ( .A1(\sra_198/n256 ), .A2(\sra_198/n231 ), .ZN(
        \sra_198/n173 ) );
  AOI221_X1 \sra_198/U57  ( .B1(\sra_198/n77 ), .B2(\sra_198/n88 ), .C1(
        \sra_198/n79 ), .C2(\sra_198/n109 ), .A(\sra_198/n217 ), .ZN(
        \sra_198/n108 ) );
  AOI221_X1 \sra_198/U56  ( .B1(\sra_198/n77 ), .B2(\sra_198/n82 ), .C1(
        \sra_198/n79 ), .C2(\sra_198/n105 ), .A(\sra_198/n217 ), .ZN(
        \sra_198/n104 ) );
  AOI221_X1 \sra_198/U55  ( .B1(\sra_198/n77 ), .B2(\sra_198/n99 ), .C1(
        \sra_198/n79 ), .C2(\sra_198/n100 ), .A(\sra_198/n217 ), .ZN(
        \sra_198/n98 ) );
  INV_X1 \sra_198/U54  ( .A(\sra_198/n93 ), .ZN(\sra_198/n228 ) );
  AOI221_X1 \sra_198/U53  ( .B1(\sra_198/n77 ), .B2(\sra_198/n92 ), .C1(
        \sra_198/n79 ), .C2(\sra_198/n228 ), .A(\sra_198/n217 ), .ZN(
        \sra_198/n91 ) );
  INV_X1 \sra_198/U52  ( .A(\sra_198/n138 ), .ZN(\sra_198/n226 ) );
  AOI221_X1 \sra_198/U51  ( .B1(\sra_198/n77 ), .B2(\sra_198/n89 ), .C1(
        \sra_198/n79 ), .C2(\sra_198/n226 ), .A(\sra_198/n217 ), .ZN(
        \sra_198/n182 ) );
  INV_X1 \sra_198/U50  ( .A(\sra_198/n126 ), .ZN(\sra_198/n225 ) );
  AOI221_X1 \sra_198/U49  ( .B1(\sra_198/n77 ), .B2(\sra_198/n166 ), .C1(
        \sra_198/n79 ), .C2(\sra_198/n225 ), .A(\sra_198/n217 ), .ZN(
        \sra_198/n172 ) );
  INV_X1 \sra_198/U48  ( .A(\sra_198/n139 ), .ZN(\sra_198/n227 ) );
  AOI221_X1 \sra_198/U47  ( .B1(\sra_198/n77 ), .B2(\sra_198/n95 ), .C1(
        \sra_198/n79 ), .C2(\sra_198/n227 ), .A(\sra_198/n217 ), .ZN(
        \sra_198/n185 ) );
  AOI221_X1 \sra_198/U46  ( .B1(\sra_198/n77 ), .B2(\sra_198/n83 ), .C1(
        \sra_198/n79 ), .C2(\sra_198/n136 ), .A(\sra_198/n217 ), .ZN(
        \sra_198/n176 ) );
  INV_X1 \sra_198/U45  ( .A(\sra_198/n87 ), .ZN(\sra_198/n229 ) );
  AOI221_X1 \sra_198/U44  ( .B1(\sra_198/n77 ), .B2(\sra_198/n86 ), .C1(
        \sra_198/n79 ), .C2(\sra_198/n229 ), .A(\sra_198/n217 ), .ZN(
        \sra_198/n85 ) );
  INV_X1 \sra_198/U43  ( .A(\sra_198/n80 ), .ZN(\sra_198/n230 ) );
  AOI221_X1 \sra_198/U42  ( .B1(\sra_198/n77 ), .B2(\sra_198/n78 ), .C1(
        \sra_198/n79 ), .C2(\sra_198/n230 ), .A(\sra_198/n217 ), .ZN(
        \sra_198/n76 ) );
  INV_X1 \sra_198/U41  ( .A(\sra_198/n140 ), .ZN(\sra_198/n223 ) );
  AOI221_X1 \sra_198/U40  ( .B1(\sra_198/n77 ), .B2(\sra_198/n102 ), .C1(
        \sra_198/n79 ), .C2(\sra_198/n223 ), .A(\sra_198/n217 ), .ZN(
        \sra_198/n192 ) );
  AOI221_X1 \sra_198/U39  ( .B1(\sra_198/n81 ), .B2(\sra_198/n95 ), .C1(
        \sra_198/n77 ), .C2(\sra_198/n96 ), .A(\sra_198/n215 ), .ZN(
        \sra_198/n170 ) );
  NAND2_X1 \sra_198/U38  ( .A1(\sra_198/n241 ), .A2(\sra_198/n239 ), .ZN(
        \sra_198/n147 ) );
  INV_X1 \sra_198/U37  ( .A(\sra_198/n146 ), .ZN(\sra_198/n238 ) );
  AOI21_X1 \sra_198/U36  ( .B1(\sra_198/n118 ), .B2(\sra_198/n142 ), .A(
        \sra_198/n150 ), .ZN(\sra_198/n153 ) );
  OAI221_X1 \sra_198/U35  ( .B1(\sra_198/n254 ), .B2(\sra_198/n146 ), .C1(
        \sra_198/n243 ), .C2(\sra_198/n147 ), .A(\sra_198/n153 ), .ZN(
        \sra_198/n109 ) );
  AOI21_X1 \sra_198/U34  ( .B1(\sra_198/n118 ), .B2(\sra_198/n242 ), .A(
        \sra_198/n150 ), .ZN(\sra_198/n151 ) );
  OAI221_X1 \sra_198/U33  ( .B1(\sra_198/n247 ), .B2(\sra_198/n146 ), .C1(
        \sra_198/n246 ), .C2(\sra_198/n147 ), .A(\sra_198/n151 ), .ZN(
        \sra_198/n105 ) );
  AOI21_X1 \sra_198/U32  ( .B1(\sra_198/n118 ), .B2(\sra_198/n149 ), .A(
        \sra_198/n150 ), .ZN(\sra_198/n148 ) );
  OAI221_X1 \sra_198/U31  ( .B1(\sra_198/n251 ), .B2(\sra_198/n146 ), .C1(
        \sra_198/n253 ), .C2(\sra_198/n147 ), .A(\sra_198/n148 ), .ZN(
        \sra_198/n100 ) );
  OAI22_X1 \sra_198/U30  ( .A1(\sra_198/n146 ), .A2(\sra_198/n253 ), .B1(
        \sra_198/n147 ), .B2(\sra_198/n252 ), .ZN(\sra_198/n165 ) );
  AOI221_X1 \sra_198/U29  ( .B1(\sra_198/n149 ), .B2(\sra_198/n119 ), .C1(
        \sra_198/n164 ), .C2(\sra_198/n118 ), .A(\sra_198/n165 ), .ZN(
        \sra_198/n132 ) );
  AOI22_X1 \sra_198/U28  ( .A1(\sra_198/n119 ), .A2(\sra_198/n242 ), .B1(
        \sra_198/n118 ), .B2(\sra_198/n141 ), .ZN(\sra_198/n167 ) );
  INV_X1 \sra_198/U27  ( .A(\sra_198/n167 ), .ZN(\sra_198/n237 ) );
  AOI221_X1 \sra_198/U26  ( .B1(\sra_198/n152 ), .B2(\sra_198/n238 ), .C1(
        \sra_198/n83 ), .C2(\sra_198/n231 ), .A(\sra_198/n237 ), .ZN(
        \sra_198/n158 ) );
  AOI21_X1 \sra_198/U25  ( .B1(\sra_198/n118 ), .B2(\sra_198/n144 ), .A(
        \sra_198/n150 ), .ZN(\sra_198/n162 ) );
  INV_X1 \sra_198/U24  ( .A(\sra_198/n162 ), .ZN(\sra_198/n236 ) );
  AOI221_X1 \sra_198/U23  ( .B1(\sra_198/n145 ), .B2(\sra_198/n238 ), .C1(
        \sra_198/n96 ), .C2(\sra_198/n231 ), .A(\sra_198/n236 ), .ZN(
        \sra_198/n117 ) );
  INV_X1 \sra_198/U22  ( .A(\sra_198/n112 ), .ZN(\sra_198/n217 ) );
  AOI221_X1 \sra_198/U21  ( .B1(\sra_198/n144 ), .B2(\sra_198/n238 ), .C1(
        \sra_198/n145 ), .C2(\sra_198/n231 ), .A(\sra_198/n240 ), .ZN(
        \sra_198/n93 ) );
  AOI221_X1 \sra_198/U20  ( .B1(\sra_198/n142 ), .B2(\sra_198/n238 ), .C1(
        \sra_198/n143 ), .C2(\sra_198/n231 ), .A(\sra_198/n240 ), .ZN(
        \sra_198/n87 ) );
  AOI221_X1 \sra_198/U19  ( .B1(\sra_198/n242 ), .B2(\sra_198/n238 ), .C1(
        \sra_198/n141 ), .C2(\sra_198/n231 ), .A(\sra_198/n240 ), .ZN(
        \sra_198/n80 ) );
  AOI221_X1 \sra_198/U18  ( .B1(\sra_198/n149 ), .B2(\sra_198/n238 ), .C1(
        \sra_198/n164 ), .C2(\sra_198/n231 ), .A(\sra_198/n240 ), .ZN(
        \sra_198/n140 ) );
  NOR2_X1 \sra_198/U17  ( .A1(\sra_198/n241 ), .A2(\sra_198/n239 ), .ZN(
        \sra_198/n119 ) );
  INV_X1 \sra_198/U16  ( .A(\sra_198/n137 ), .ZN(\sra_198/n216 ) );
  NOR2_X1 \sra_198/U15  ( .A1(\sra_198/n216 ), .A2(\sra_198/n146 ), .ZN(
        \sra_198/n77 ) );
  INV_X1 \sra_198/U14  ( .A(\sra_198/n109 ), .ZN(\sra_198/n234 ) );
  INV_X1 \sra_198/U13  ( .A(\sra_198/n105 ), .ZN(\sra_198/n233 ) );
  INV_X1 \sra_198/U8  ( .A(\sra_198/n100 ), .ZN(\sra_198/n232 ) );
  INV_X1 \sra_198/U7  ( .A(\sra_198/n169 ), .ZN(\sra_198/n214 ) );
  INV_X1 \sra_198/U6  ( .A(\sra_198/n147 ), .ZN(\sra_198/n231 ) );
  NOR2_X1 \sra_198/U5  ( .A1(\sra_198/n216 ), .A2(\sra_198/n147 ), .ZN(
        \sra_198/n81 ) );
  NOR2_X1 \sra_198/U4  ( .A1(\sra_198/n218 ), .A2(ct_1[5]), .ZN(\sra_198/n79 )
         );
  NOR2_X1 \sra_198/U3  ( .A1(\sra_198/n239 ), .A2(ct_1[2]), .ZN(\sra_198/n118 ) );
  MUX2_X1 \sra_198/U226  ( .A(\sra_198/n202 ), .B(\sra_198/n235 ), .S(ct_1[4]), 
        .Z(\sra_198/n201 ) );
  MUX2_X1 \sra_198/U206  ( .A(PR_1[31]), .B(PR_1[30]), .S(\sra_198/n124 ), .Z(
        \sra_198/n149 ) );
  MUX2_X1 \sra_198/U142  ( .A(\sra_198/n157 ), .B(\sra_198/n158 ), .S(ct_1[4]), 
        .Z(\sra_198/n156 ) );
  MUX2_X1 \sra_198/U115  ( .A(\sra_198/n131 ), .B(\sra_198/n132 ), .S(ct_1[4]), 
        .Z(\sra_198/n130 ) );
  MUX2_X1 \sra_198/U106  ( .A(\sra_198/n116 ), .B(\sra_198/n117 ), .S(ct_1[4]), 
        .Z(\sra_198/n115 ) );
  NOR2_X4 \sra_198/U12  ( .A1(ct_1[0]), .A2(ct_1[1]), .ZN(\sra_198/n124 ) );
  NOR2_X4 \sra_198/U11  ( .A1(\sra_198/n255 ), .A2(ct_1[1]), .ZN(
        \sra_198/n123 ) );
  NAND2_X2 \sra_198/U10  ( .A1(ct_1[1]), .A2(\sra_198/n255 ), .ZN(
        \sra_198/n120 ) );
  NAND2_X2 \sra_198/U9  ( .A1(ct_1[1]), .A2(ct_1[0]), .ZN(\sra_198/n121 ) );
  INV_X1 \add_35/U1  ( .A(q[0]), .ZN(qp1[0]) );
  XOR2_X1 \add_35/U2  ( .A(\add_35/carry [30]), .B(q[30]), .Z(qp1[30]) );
  HA_X1 \add_35/U1_1_1  ( .A(q[1]), .B(q[0]), .CO(\add_35/carry [2]), .S(
        qp1[1]) );
  HA_X1 \add_35/U1_1_2  ( .A(q[2]), .B(\add_35/carry [2]), .CO(
        \add_35/carry [3]), .S(qp1[2]) );
  HA_X1 \add_35/U1_1_3  ( .A(q[3]), .B(\add_35/carry [3]), .CO(
        \add_35/carry [4]), .S(qp1[3]) );
  HA_X1 \add_35/U1_1_4  ( .A(q[4]), .B(\add_35/carry [4]), .CO(
        \add_35/carry [5]), .S(qp1[4]) );
  HA_X1 \add_35/U1_1_5  ( .A(q[5]), .B(\add_35/carry [5]), .CO(
        \add_35/carry [6]), .S(qp1[5]) );
  HA_X1 \add_35/U1_1_6  ( .A(q[6]), .B(\add_35/carry [6]), .CO(
        \add_35/carry [7]), .S(qp1[6]) );
  HA_X1 \add_35/U1_1_7  ( .A(q[7]), .B(\add_35/carry [7]), .CO(
        \add_35/carry [8]), .S(qp1[7]) );
  HA_X1 \add_35/U1_1_8  ( .A(q[8]), .B(\add_35/carry [8]), .CO(
        \add_35/carry [9]), .S(qp1[8]) );
  HA_X1 \add_35/U1_1_9  ( .A(q[9]), .B(\add_35/carry [9]), .CO(
        \add_35/carry [10]), .S(qp1[9]) );
  HA_X1 \add_35/U1_1_10  ( .A(q[10]), .B(\add_35/carry [10]), .CO(
        \add_35/carry [11]), .S(qp1[10]) );
  HA_X1 \add_35/U1_1_11  ( .A(q[11]), .B(\add_35/carry [11]), .CO(
        \add_35/carry [12]), .S(qp1[11]) );
  HA_X1 \add_35/U1_1_12  ( .A(q[12]), .B(\add_35/carry [12]), .CO(
        \add_35/carry [13]), .S(qp1[12]) );
  HA_X1 \add_35/U1_1_13  ( .A(q[13]), .B(\add_35/carry [13]), .CO(
        \add_35/carry [14]), .S(qp1[13]) );
  HA_X1 \add_35/U1_1_14  ( .A(q[14]), .B(\add_35/carry [14]), .CO(
        \add_35/carry [15]), .S(qp1[14]) );
  HA_X1 \add_35/U1_1_15  ( .A(q[15]), .B(\add_35/carry [15]), .CO(
        \add_35/carry [16]), .S(qp1[15]) );
  HA_X1 \add_35/U1_1_16  ( .A(q[16]), .B(\add_35/carry [16]), .CO(
        \add_35/carry [17]), .S(qp1[16]) );
  HA_X1 \add_35/U1_1_17  ( .A(q[17]), .B(\add_35/carry [17]), .CO(
        \add_35/carry [18]), .S(qp1[17]) );
  HA_X1 \add_35/U1_1_18  ( .A(q[18]), .B(\add_35/carry [18]), .CO(
        \add_35/carry [19]), .S(qp1[18]) );
  HA_X1 \add_35/U1_1_19  ( .A(q[19]), .B(\add_35/carry [19]), .CO(
        \add_35/carry [20]), .S(qp1[19]) );
  HA_X1 \add_35/U1_1_20  ( .A(q[20]), .B(\add_35/carry [20]), .CO(
        \add_35/carry [21]), .S(qp1[20]) );
  HA_X1 \add_35/U1_1_21  ( .A(q[21]), .B(\add_35/carry [21]), .CO(
        \add_35/carry [22]), .S(qp1[21]) );
  HA_X1 \add_35/U1_1_22  ( .A(q[22]), .B(\add_35/carry [22]), .CO(
        \add_35/carry [23]), .S(qp1[22]) );
  HA_X1 \add_35/U1_1_23  ( .A(q[23]), .B(\add_35/carry [23]), .CO(
        \add_35/carry [24]), .S(qp1[23]) );
  HA_X1 \add_35/U1_1_24  ( .A(q[24]), .B(\add_35/carry [24]), .CO(
        \add_35/carry [25]), .S(qp1[24]) );
  HA_X1 \add_35/U1_1_25  ( .A(q[25]), .B(\add_35/carry [25]), .CO(
        \add_35/carry [26]), .S(qp1[25]) );
  HA_X1 \add_35/U1_1_26  ( .A(q[26]), .B(\add_35/carry [26]), .CO(
        \add_35/carry [27]), .S(qp1[26]) );
  HA_X1 \add_35/U1_1_27  ( .A(q[27]), .B(\add_35/carry [27]), .CO(
        \add_35/carry [28]), .S(qp1[27]) );
  HA_X1 \add_35/U1_1_28  ( .A(q[28]), .B(\add_35/carry [28]), .CO(
        \add_35/carry [29]), .S(qp1[28]) );
  HA_X1 \add_35/U1_1_29  ( .A(q[29]), .B(\add_35/carry [29]), .CO(
        \add_35/carry [30]), .S(qp1[29]) );
  INV_X1 \add_34/U1  ( .A(nq[0]), .ZN(nqp1[0]) );
  XOR2_X1 \add_34/U2  ( .A(\add_34/carry [30]), .B(nq[30]), .Z(nqp1[30]) );
  HA_X1 \add_34/U1_1_1  ( .A(nq[1]), .B(nq[0]), .CO(\add_34/carry [2]), .S(
        nqp1[1]) );
  HA_X1 \add_34/U1_1_2  ( .A(nq[2]), .B(\add_34/carry [2]), .CO(
        \add_34/carry [3]), .S(nqp1[2]) );
  HA_X1 \add_34/U1_1_3  ( .A(nq[3]), .B(\add_34/carry [3]), .CO(
        \add_34/carry [4]), .S(nqp1[3]) );
  HA_X1 \add_34/U1_1_4  ( .A(nq[4]), .B(\add_34/carry [4]), .CO(
        \add_34/carry [5]), .S(nqp1[4]) );
  HA_X1 \add_34/U1_1_5  ( .A(nq[5]), .B(\add_34/carry [5]), .CO(
        \add_34/carry [6]), .S(nqp1[5]) );
  HA_X1 \add_34/U1_1_6  ( .A(nq[6]), .B(\add_34/carry [6]), .CO(
        \add_34/carry [7]), .S(nqp1[6]) );
  HA_X1 \add_34/U1_1_7  ( .A(nq[7]), .B(\add_34/carry [7]), .CO(
        \add_34/carry [8]), .S(nqp1[7]) );
  HA_X1 \add_34/U1_1_8  ( .A(nq[8]), .B(\add_34/carry [8]), .CO(
        \add_34/carry [9]), .S(nqp1[8]) );
  HA_X1 \add_34/U1_1_9  ( .A(nq[9]), .B(\add_34/carry [9]), .CO(
        \add_34/carry [10]), .S(nqp1[9]) );
  HA_X1 \add_34/U1_1_10  ( .A(nq[10]), .B(\add_34/carry [10]), .CO(
        \add_34/carry [11]), .S(nqp1[10]) );
  HA_X1 \add_34/U1_1_11  ( .A(nq[11]), .B(\add_34/carry [11]), .CO(
        \add_34/carry [12]), .S(nqp1[11]) );
  HA_X1 \add_34/U1_1_12  ( .A(nq[12]), .B(\add_34/carry [12]), .CO(
        \add_34/carry [13]), .S(nqp1[12]) );
  HA_X1 \add_34/U1_1_13  ( .A(nq[13]), .B(\add_34/carry [13]), .CO(
        \add_34/carry [14]), .S(nqp1[13]) );
  HA_X1 \add_34/U1_1_14  ( .A(nq[14]), .B(\add_34/carry [14]), .CO(
        \add_34/carry [15]), .S(nqp1[14]) );
  HA_X1 \add_34/U1_1_15  ( .A(nq[15]), .B(\add_34/carry [15]), .CO(
        \add_34/carry [16]), .S(nqp1[15]) );
  HA_X1 \add_34/U1_1_16  ( .A(nq[16]), .B(\add_34/carry [16]), .CO(
        \add_34/carry [17]), .S(nqp1[16]) );
  HA_X1 \add_34/U1_1_17  ( .A(nq[17]), .B(\add_34/carry [17]), .CO(
        \add_34/carry [18]), .S(nqp1[17]) );
  HA_X1 \add_34/U1_1_18  ( .A(nq[18]), .B(\add_34/carry [18]), .CO(
        \add_34/carry [19]), .S(nqp1[18]) );
  HA_X1 \add_34/U1_1_19  ( .A(nq[19]), .B(\add_34/carry [19]), .CO(
        \add_34/carry [20]), .S(nqp1[19]) );
  HA_X1 \add_34/U1_1_20  ( .A(nq[20]), .B(\add_34/carry [20]), .CO(
        \add_34/carry [21]), .S(nqp1[20]) );
  HA_X1 \add_34/U1_1_21  ( .A(nq[21]), .B(\add_34/carry [21]), .CO(
        \add_34/carry [22]), .S(nqp1[21]) );
  HA_X1 \add_34/U1_1_22  ( .A(nq[22]), .B(\add_34/carry [22]), .CO(
        \add_34/carry [23]), .S(nqp1[22]) );
  HA_X1 \add_34/U1_1_23  ( .A(nq[23]), .B(\add_34/carry [23]), .CO(
        \add_34/carry [24]), .S(nqp1[23]) );
  HA_X1 \add_34/U1_1_24  ( .A(nq[24]), .B(\add_34/carry [24]), .CO(
        \add_34/carry [25]), .S(nqp1[24]) );
  HA_X1 \add_34/U1_1_25  ( .A(nq[25]), .B(\add_34/carry [25]), .CO(
        \add_34/carry [26]), .S(nqp1[25]) );
  HA_X1 \add_34/U1_1_26  ( .A(nq[26]), .B(\add_34/carry [26]), .CO(
        \add_34/carry [27]), .S(nqp1[26]) );
  HA_X1 \add_34/U1_1_27  ( .A(nq[27]), .B(\add_34/carry [27]), .CO(
        \add_34/carry [28]), .S(nqp1[27]) );
  HA_X1 \add_34/U1_1_28  ( .A(nq[28]), .B(\add_34/carry [28]), .CO(
        \add_34/carry [29]), .S(nqp1[28]) );
  HA_X1 \add_34/U1_1_29  ( .A(nq[29]), .B(\add_34/carry [29]), .CO(
        \add_34/carry [30]), .S(nqp1[29]) );
endmodule

